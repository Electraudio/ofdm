��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��p&%CX�WD�m�;���2��A�Z+k��H����+a��|O��g�o�c�l��w&Y)Lk�֯�#\��h�=x�PA'��N��i.�l��Nb�H��x?e��֍o���
�B���;�u|Q�6:��0��w����)Pغd(F8݆p����� p��賘4/�]?���=pS��;WƵa�*����S-3�kH�~h�i*�4[E�Xi$k�;�;��s��$:ٜٛ�,��S{y��(ХO����Q�r*��L
�a=gj�]��*�t��R�	�P_�p���j���o;��p�6ВT��������m2͑_��c� g�0���x��$���b�ݭ?Ti���3׮�"TԜL�zi�UZ�%�mAJ\��5�����4�T3����I���a�@��t�{-\�z�L���E�� m7'���n=���Q\C?�@$G�f
C����I�����jaw�}�1@�+�fH'�.<b�ĵo$@X�=CB[j�7��*y�+X�fj�}�VQ��
��㟄S�����sxh�Xq�3��n��r��IȣF�	���
��}	P�$����1Z�ǚ"RU�Ǡ2^��y�d�]��t��ڞߪ��2op��W
T���<V�'����_=Uf\^�	��/� �
i��/L-��Wb��2���>}L������>�D��H����V?��7�Ĭ��M��e�A�K�ѧOY�j��P�gZQ�=Y>L�O�yM+�h�q�t��m"�T�6i�F�X�F�uT+���t6�Snn2D�O5	>(P��u8:����X�������v}���x�3�����O�����m�Ɂ~HE1v�M���n*t�IOn}
:��A���]Ҩ�qB0��JV�rS-TU�k>
�_%ه�(;�μ-�}M�EO8�a�sr����EÑcb��Agx��i�!�I����N�W?�
����/BP���ڥ!�`���K$�2�ث�zbWTJՓ�����AI��'.�:��i)��b��h�X�9o�]}>���\��`��m-~�>id�,X:@��R���4�8{m��߾�Z�0S�N
�������� 8p���T��d��١��LǶD�j	��f�E+喨W��T�*�ާ�7�-����9w��Kt&��˽��=|A*�G�
C��9u�0"sqg?u���s�D:Ò������P��)�Ƃ]2Q��גKA�ã�� sV�w�����^�<vka��oAً۟R��4����-ɶ�<b)\7�}�:��;���):Ħ
�n�s��>�? A76G��la3}�r�ҙo;��V�U	�h�b�~疨�?R�X�� ��t�6l�U�M?0`�)ʼ)L����z%�2��-0$5#�d��}[=O�g�}��4p����v����q��)�n�-bh% ��@Lrj;�)����`D@�DvR�6�I[�*���}�M�� ���yc��;�z	rNNW�	1��J���:�x�?]���e���Ծ���<�̧D���6֎�IX�'���+a�ֈq~1��&]ߞ�y�Ld�����B`�n�S/s>���䨖}fu<���(1��8�f��J�;�g4;)f�@wMP��Y�Q����7tCT|ʰ���ȅ��8e�9�Ŏt:������D�1T��;���FW%t w�و��q:N��%ƹ(\�b�U��:U}H�*�՜�9��>�`Y>���^�$�e��^��I�µ
��M�wҚ^��[��MS���q�+�f^���sK	�Z�Dt��;�6����ow&\Q"�0��|�Z~����I���ޮ�L�4�.�s$����`��$ �ş��{�Z/'Sl1c]��!Du�^�2ͦ�/��\�� ����Q��C$����(1h�1��:��O�|\EF��m�i���&}�$�b�δ���m�{m#h�Y������7��k��j��}�J�*��+���f��s��U)�W;YU�T��Z��5��fh_���܂ZTo���]RF���2�D<Ⱦ.+�0KhjY4�Zt7��m��3@�6�&K��@�@B��Mg
u���S��}�T�d%iy�q��9ȗ�EM�����lM�%1g�GXX��!��]ԡ���@6f�#�gK�EW�P���y-�l,<ƷΨcȜa��Lt��=�I�%����ٞ�5Sn'�03o��:�.����}*M��� VYG��z�٪s̀�p����[�CH��7�ǥH�	kO7�E��#�Z�=H�Cȕ���dz��y�ᗙ�S��hU����+�ꀀ
�n�uT e��<��P����Ҁc���!#.�?�T$wK�-tq�.�K�LZO�������N��Cf�X����"��Gva}2Y�tQ2�ҸP���?���M��l���}s.�h������'y�w�Z$쫐��� ��~+�־�9dh(�|�L.����=���zyd�.W��\ Rh�k $E�U��-\�ܥ���zj�!��Vr�a	˾�O �r�!�Q��*�M/��m���ߥ��@���W���j��,�L[��I�8��=_uR�)_�?�I8�1-K�p�t's���Ш�ܛ��;_���Bu���)"j�B��|��#��a�� /�;4=�ߥ��8s1��ѝTD;,K9 w�-�^�&�)Ha��P�GBP�1��GhjX�R��ak��$4��Ǐܛ%<L\��پ�+z�r� ���Z��F�l�	��4ʟU�P���Ur�5�	��r�ަ�e�T�):�Io��a�®�p��XDrmI��il~�ET��d_�j�]>Ue�<-9�6��JvA�b��oS��c�tm&�����k�-��cN��P�ȕ�V��4�Q~=S�=�-Ui�? dD�꨾k�$�4��Nu�"��O+m� !��d�AϘ�i��w.��Yv�J�M�_���Q�҇��36��Kxǭ+?R{5���b���������
���Y��q����r�k����M���*�	E��"������6�τ���T�B���9���V+���/��>K������S����53 wvP�`���C:[�xd痿}� � ��9��R��|������F�csz;:���X�':(�|�J�}�H�C���o[�3ηS-���Բ�e�Y?M&Y5p�6��G!0s$0��Y9��>�o9�ek=�P�ܢ�ټ|���{�l�