��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`h9�_�p^Ku5���>c�r��.���g�~"ͧ�mj��A��j��(	e1�K�߽ώ�q�O"ð����u��Ǜ^֢��p��TI�1��m��	�@g��1��Ii����Sϔ���P��Be�r/�8׹I^�w$����iv\#	��H�܆ej�i�_��O)�I���pGǘ�ﴵh����H��d�&��?~�d�)J�w��QP`���z�a�x��&F֧���7�q����!�%h֗hV^:w���R���ֆL��#s�H4BԅZ ���)jDN�r��g�n������&�j ʱEy��p�Er�mƨ��Q5A%-^sU�9:͈��㬟4��b����5��:��E�NX� $�x(����:�ۉ�p���}
�����=O����n�d��/R
,�ۖ�P� }'nN]Y��w���*�b��b�Û�7�
�g����I�l�~9�����}�1�:jp|���b@��V�À����ޢ 1'�ɻ��{��Ȇ��
��P`���S\25�๲Y�؈�&ez<�Mxr.�ӭ*��Z����&�B{;�F�_�;�Q�c&�/�W!"�����[8��%�����P�2��m�r&�U�f�J?�����u]m���v�Y8�}t��c6�`��iL6��Tr��V��IzqLMQ�a)�c����n.�:\w����	��kP�A��kA���a��MA�*��;�&�y�Kpc��%{�\��`]ޑjLe���]��y߼����o6f;S"Z���]KG�Q�6�ݧ��y*g o�[O��.3I���x@N��9�8 gh���ww
)�ا�.q�Lv��'�9ݻ����UV�u��^٨:�}���|ӻC ���4��	k�r0����dc�x�"���)�W�;�n�,��L�q�_��EѾ��7��6��J韕��\���zqY��FnD��:�4DI����q�l ����X�T��k�i��&��*�'�	fA}G�%>�9��yO,Er�8��ҧ=�x���Dz�MܨRA��a]�zԜ��bJF9����|�?\CE���v���ՐS��^����������`��L6��hU�=brSV�j	44�L�����m��'�E��!� ��F�!��2��!D�Z"�_�3�ґ�����nQ,�:�G�.52��0T������H�Q�R4 3��U �--�"�����C�e����k�	E��aV�P����s��]Qp���Y��=��>D|�W*�/�[�=/��G���q�m�7�u�\����Zz�k,��h��l�O��!ʹ�v��wª1�'�kS��6�7~� %�"&u
�n-7�MQU�*B�ьQ�zD=�t�����]���^ơV�����k�d��g�ӆ!�*}�xSr�qΈc��Yըs���G*��q/� �s���.�� �M0n����ѓx�kML���j�X����dr�֛�J��������ݵ�!���/�p�
܂AR.�2�"��x�z��
j�oR��P��[�|�@#:y	���z5
`�����4e̍h�&f~8��|*;7�Ŵ���;,�;����c�Ik�F�}��Hu'�GE�s�����P��V��d|�]�ѧw��-+�VS�3?EŇ��ֱ;D"Q@M�p�;�ѷ�Ex/uV&��b+��N�61ǆͧ��$!�U|Җ�SژY�Sr����{�$Q�6�Ȇ�E�g���?�|�kU`z�Б��/�&�;��%4�HCvu�8$�|9�]=8��y"�4''�.i{��;ha���_	}f��0���҈�\��*�Bf �71|ZSc(�­�S����@�5�C8��Hs�lR��|��5)!y�_8�,Yͩ¾�M���	%bP�,�B���U��J��*�D�4˛X��6%}@��p�E�횤��'b����v����(��wKG}��AݰQ����gW9ꜘ�#��S������ܼ�]�X��^����חS�J����ˡ��M��;���h�(�՟�䮺5��]`cs�*r~e��8s6}A�V�ϓ�0���gQ�6��UNW �ߦE��s ����ˋ� W��=����`�>�	9�ت��D&m�U���8f,
��=�˙e'S����1<C̾7@�Kq`'G�(w������t��7W8:�8�����?�zT�XY�3:D{��ps/�(�?u�	��.e����->����@yy]�0G��X)���ۥ�~5��.�3�t
=ɹ�J�?#���YӴJ-��k�ʰ�k~bS�鈍f��|�d��^��(e���{j�翮]�����HS�9���|q��HB�z��6�Az�G�YP<��}P��L#Nt�Vp�Y�_?���3�	4)�ʷ�D�@��~%&�]�eR�}h�bY	<��i'����ŔR�������:V�@�"% m�ku�X�r���f9����u�0ה~��l�#��W�q.�@G���us�숇�% �g��߸�����ѾU~A���6+�d������u��\iwr��I��y�"�|����9��k�[�Y^�IZՕ^���!Q'&�C	O�n�7As�?�ю,^S��0�,D���O߹��^���
�?�'ځ������
�����H#��七pI>R%Ls�V�*ޏw�����A�ŇU?�N{!y����a}X�1q���W���>��>�b��Q�:aO⩐�zW.O�R[�f2�����孈-�=N�.�RmEE����^r�a[f��&#�m\q�`�e�Bf��+_����m'�b����,���mf)y���Li�R[�!(I�TF�c^�!��'N�����^��L��7��|ŰpiME.�e�L }�9��ю/p�͍��p��2(�+��� �P6->��I �i�I��3|��QB��a�
\��d�V�[��t#E�G!�zi��W
?�:�P�фZ�˚����>��d����̓9Um�_Q0���4"��H��s=��W�D.��z��ϖ����EɜvԠ�4������K%9�u��띵j]�
 uxu�"��F�Iy]��3�0�ȫک:,�e5%�g3=;T��=��m�^Rt��.�M�����4�.��3�&SP�d׊(E@��9��1 ���ʍ]���	��7�Ũ�Y� 2�Q"��9;��r����W��ւ�!>8�&�j.<�&{���:ɹ2��\���1+���'IAuf�� �Z�N�ɻ�`n	��O�g~~n�@Y���Ö��^�B�ܨ=^��s���4��?�F�����@>v�����M�B���`����N����$�&�l�����D(v��K�\�p�z�@��tz��,nkM��I��8��t'���Rf�0�ǁ��C$�����q���M8p��~]D��)��L@?7>����ީ�Ӝ=�Pu��ޣ�k����r�9p�Y��=�:���̠m|�����27cL�4ӹ#�~�;��v�Y,/} �������L b����\��n����(��wg��/
=٠���Gmxa2'$���'�_�7V�/rI�����t�� ��u(����
4'�>_,��Ԡ�$��Tz�^��ň�=�b�
�-��x"��xh�q���Oύڈ�V+|h@�Y����������#~a�T��YڇЯ�����ý��ժ]ԀN+ɮ��K��_�ݽ�KރϏ,}ʀ���`;���W-^z�p<����'#��1����fL��6�_�.�C����	��!�DJ �b���>�v�1���y����/-��]F͆�P�?R��xE_��m�䋭���z��	('b0f�;f���M��S$&��i�0�����u�m���<�L'6�#�Ɠ�������������r�ӍP�x�m�:ʋZH���%U�D�c�eÌ^v�c_;{�J�T�$\���/U~�D�?���B#���~LVW8,�18�K�X��%������nI�$)7�C�MeFBX��3<�GJ����F�#b�$��b��^���e=�R���Б��\�9���-��4�����ZĊ�����-A�}N��ҍq<�I{XX��z�N���l
������l�ܷ��&\�����qC.`Lտi�54/�N�E��&�nڗ�JQi��ҭ'��u�5UGN���	�%ܻ����*��ys���#^�7����1�`S��3<��a�X/�����Di�)�&��HO���@)�
�����s-p� ��(=�zA��oc��?)��}D]����wO��vV�� 7�skVƷEU{��XQ~]�߮Ҳ���:��H��4&_">�ҧY�.�Q?�{�/;E�$�kT�E��w�]�[ ��Q���=��������T��_��UM.?����o�~�A��,���Zu�_���j��ȴq�Uh�cȀ(�[7$�g����)�hc9�|� �n��U��mBpy�Xyq�ZX^�۔�����փT�K����b�sp����Qض���/�b�?�'�!I=��t`;	�����<a��=�����\��4[��*��(C�V� [�(�\���?mޠ���	�w)�>G��yRi��bU�O�}�P$�Z�`6b���hF��^��	��	Xޗ��?�EE}��n:J���o��!��p<�S��NE-}��i���K{ہ��KY\-V�5k��C��!��Փn��M�͑Z��<�>�h�Щ0����|TPϊ �fz.M�a۫)JTG-ͭl�$���k���~��?V��y%��L8f$��� Ҕ�2�����ϕ>�q�bA�g�UWS�XW/��a�"�{��w�!�v���@��̽v��˻�U	jdbGi��`}U���H-��~�;�xj�$�;��7�9��Y�MA�5'e�`k�N�s�����-���y����ⴽs�Iͱ�����Y곅�O9��X���D�b�j��`ĭ��5�~C�|�y2Z�b�]�#t�b�{��jtm/P��Ax�B�?�����-�H'�P���죣t�s���@N��a����I��J��?؀ù��@�+1�*�!Z�T�(z�R�C0%�eV:*�l/��[բ6)c�x�@r��ւ0�o)s.����꿩��O`xFC���wW�pw�6����>��X��e�����xPQ�ߦ5��Nҷ�D����t�ct6�8�7ճٿE�@��a�m���":If��	��u�_@�r���D�2�B-.֭ �;nJya:<�����-��HwД
�PV�	�[�'B�7]'��
d���L<vhh�bA3���/���:�M1�<���
��ciN-|z�v�N/��ýu�(��Hd8��+^7_�iI��z���s��N]������T	�}u�C����%ebT�k\U�2��-�B���^8�bGTB�<w�G_�Ə�B�A��غ��G	��M*,{/f��f�g���������U�Ƃ�mQn����B�2$�\���n�P/q�=r���ܾzM��提���͔� �_�l\;0�g�L-�z?���']b(Ǫe�֟�+����\��ɼ�і�R�S	@Y�;c���������-���z��W{��&@�"����b�T��׊�r���n2ѷ�c�QJ���`��W��������R1%{	|����F���	I����O�Y�	��L^����潄�i[w�P��8Nyr�f�R�o��8Gփ����mL��O�߽�,[Y��@�4^+u����c�5�[
��>n���5τ��Z�gK��7�hV74J��ޜ}d�~�ooZ��o�����7jBдb�k���r��d82M�������WaLQ5��L���T�O?�r`�޻N�nVQ���e<�l�����"�+�������~��
��i�&v�z\���^+_�Ĺ���:�?rC��Z^oL<_�sDCO��u=�ė�([��63��%yg#rVs_o�%y'�ޓE~?V�q�����4�6Vɲ��X� y!�|��х��3֒�W����k��#�	��5Ԍ�"zI�V��i��q�C~&uR��I��	��8H*+h�)~8������Q��pd�YJ>z,��I,!5'p��5ܷP.-D��^���¾�Ľ���0����������䰆�"N�ُlE�!w)�I6Z`\�R�; S��NB��{FIg�MxF�mV��#�����r�N"ό>��������K�`�Vye^ob1K��έ�{�ݭ&���*�HUw�٬itgy�Ŏ����a�0�B�IW5�����؂���m�����S�K/�P9�ې��1��q	Ӷ�W�:�L�j)L�I��'�"��Ӱqz�=O&}�1
,���	ܩ���b<e!R9Z�5�����˦��,phh��4��p}"Bj�]�r�t˓��G$Wn^4���~���J�����[���v'2S*sbN%n��bK⃊"&�0�M�|��T��pK��������s���K7��r��U�¸���&	��+�K�nʨ�AE��S��S�J�/�f4>����!�)���H��5��ˎFs!8A�qC���jf���Ŵ�Qi���v��(l���\(�����{�3�#�����F. HY��(� ���� ���i���K�ں���h��	�������sB��Y�X���*K����&	9�X0<��<՟!�a)昤A��)��r_S�J�N�� �\,{>�F��-	$�����_6�;�����t]��I�Ov��(���ʁ])�)م��=����� עW4ۧ&A�Ikt:y���+�_"L�%�?gG�Z���~�}����� �ān��w���C��l��Y��8�G�Ժ���f��y~���NV����,v6Њo�Qf')G��Z1��tf ��o�Tq���p�:]�oC�S�t�*�g'�R��`.H�u"�"�*�7��-6;��FQ��e0��	��5PKwi�ş�@��-�_�p����d�h�TUwܗj����<��s���(��A*Hl��r��o��u���t30ʑ!���9�0M�L��^p��G�65v���S�װ��A��&zmZMhR�"-'F���^��{KN�ۣF�Gud%�i}��3�I���!��l-�W��r��c��}�����H|�)����?�ҷ�͜.��l�y*��`<U���>-Z����l<�#*�M�O��S�B�o�O㊝A\�=+$�Ђ��oG��ӈ7�>��l�=/���wj����y��	B�A��	��54��9�ܱ�����_�-F� Obǫ�;��I�Z 5���A��h�=9����1�;G��>���M�'�3��	�chP�
d��z���T�8A�R��L*ù����ɞ���l�� i��M��͟�[�?W����U��a1hؠ�a̵�a+�@�c�+�J1�ˌ#����T)5��?=�3\��s��Tq�ٗ(>Q�5Vh$]�][~R�ݠǄ�	� ��i��96*��D��^Q����`n��xS�s~��_�#���iT��W�]�J�ua,����I�Jq]aO%(QeI癑XT3�q#R�1�˘M�v	����~�5l,+QO��&h�Za�*���Fh��0�8��i�j8�V13�󉲸t���,r�du�{��}�u���{{�bk���s��T��6U }i/��p����sV;3��"kY��)�֎���P��o{ҙ�I��H��q��W���XY���Z�%���?�%)K'�M�$�a������){�X�c�>⬄{̲��9���f�jh5я�"Z��3���5ΐ�3aE��O2Pp[��&	'�u���4�頧�.Ej"�s��4��&lk���ã�R����<��H��R�V˞i$ ~�_���t�>�GM=(��»:����Ut��a�!;�V
 {���~J�~j6��6[�_첿�u�6sA��7�t�e�"�sy��1z�c�Ǒ�&�X[+��k8��IK��:!���n���/]������/v�`�Ρ!����k䂠#8L�޾wG�Pg휘�zO�:Xr�7y�+�*MS�zRudq3��K�IO��:�P��K�x���V<evd��W��suqH~_qџ:K��W�'�@Rq����Bvp������$Hh2��U-]a3��~�HǍ܏����Q��[�0�ө�����ˏϽ�u%V�H��?�4m�~�
�7��;�F�h�`�����ڷ�$J&*N�H���"�~"��@��$V?�:��2�ğd�ʦځ/��?�I����WU��E<J1�3]�1���r���S,���{O���9�&y�Or�E�39���[0���K$�d<�	�ˮɐ�S��"��Zr�
�i+�=s�*���6}ޛ#O��拴¢}�/�`Ǽ��İ3�py3�
,W*~.NW�T�nfI<%:�����^'����(l��w1¾�R6�	��f��5)�1MTey���8�?]}o7R���ѣp<y��B8MI\�e�����ְ��oa��{r�/Ci4�&��J�}J�}B[�I����k����9�4������.�گ`B�T���VsԔ���j�5SH�[��Rw�΍��K�B���ԃۯWM��0Ο�q�L\�	�����B�q�����ϸ�ˮ�9Z��EX���C\�/�Gټ܈5a����R8 "XQ%B�G!(���L6�<��9c��s���R� )1����i��:�|����(���CC�+d�T�~z;�������<���.�T��lN�4zd� <vWt`ղVp^v���Q�$�J+�o�V:��ㄌ����*�c�tF3(lW,@c�-'M��)8��!���Y2����,�2��н��	�/ؕC����q��(�g�:�:ry3I��}l�MwVqۼ�}s4��?W`�ٛ�BWˏ�t���e�*���5��BQ�Μ�>*� v"�6�z�u�z!��C�eZt/�����Ιt����(�q\���GM�q�!6;[�?�<O��pҒ�w#	V��� ��l^��^����UI�׈/�2#�}���+��u����\o}�:�}�bz�؟Ƥ�Ȃ���^o/#���2�pK|,`�\�A`(��t�`W»bq�"s�Ȋ�����)���>y�R�B#5]���HO2�Fv��"j��!*B���v��~]t�����6��=��Sݲ�`(�֚���]V��:��I�&G0�$�V�>XV���	4>+(���Ix*�V[�7�HD=>��ƫ,a�C���4`w��jZ��{�}��&w�h;�����}�w,�n�ѭL����Ձ���H�W������\�2���YQ��;2�B�Zŝ���{�[�#Nŕ���pp�~����
�kU��;�`���us���!�c�Ԅ۳��_Y"i!L/�j,�7PH|�{Y�T�BA7AtO� 2Ϟ�#�A=`�K�R����e�se�ݳ�ԬTG�ʯ��-X��2���X�"ml�(��yF�����v����4P�b��v�.���i����>wq��f{����~��CGP��a����r��X�7%��Ñ^0����n<��?�!C�;
��G;#"H��4���kN��2 aX�����T�V�~v�Q��a�7[�0|+D�(L��� *��^����7��jǝ�7%�hW�E�N��PL���݋@J��1)���B%�� ���J��8�#@�>.�g`��Iۇ�'���q8si*P	�LkK
��4Ql`d(�酣+�@���tK5�G���.�<���r��į)��H4�^e1��`ш��V�F��b8fҺ�UIT���,2X�H�����	d�0f��ߘ�Wtg��)G"�`?x!�5�B��,��MI���Ӂ�R���7WdC�+oW�,�xex���8�������º:S
e/RA�*��/X:��R -}tW����,5����)z��0؄h�G��@DɁn�����֪Sv�-B �OUD�����Sr��lu�Cs�Z����Q����&^��W��ɻt���d )�8�]�`]���}���y�~	RBD�A����r;��'��:)�bZ{��LH���&��>�6�x�L)�լ'���&^:Վ�q����Q��������۽])}*����N��~P˶��a�Ųj�i��ӊ����g��v�<$�T|P����`�1��1��m���N�q׎1�[�S?	��
g�y��o�
�r�@�G˄�A� ���s�0��_�y������WvGSTڦoL��B��ļ���Sa�������%��4}p�!�^�x�A�u;ӆ��i��3Yc3��>)BS�$҃��t�o�3~�REѴ�H]�h��DJ����0�c���
���9��v�WY�K�	)Y)P�Z9�ԑ�E3:ǹzU~x)���~ZqeJ*�^�͈�dDF��r��g�l�A������:ધT�E���l.�-�b�	��-%�o����|��߼P�|�LxD�y_o��i�՚X͛�(B�+�:[m܋k~�߭ �+`��iL�Y������!���4��f��%�b x+���w�m�1��Ɖ871�&C~�3[�}���׮��,�`�A�ıg�Ϫ��vpujV�:��\D���s�s|9���ƘzF���u~#�X�l�M��v��=���6�1���٠�C�{�I�x����l�<�^i��6~�����!��_�Q��v�I�2@�c�D%��3T��\���#s�r~?R� ����b2yU�/d�|���%\�L���x�mD�Ǟ����8�~����|ѵ�NY��V*8b	������{��m�h�a+�!BUn�{A��i]Z��AJ�Ӻ��C�$��9���^��4����2z��fg �/G�*k���"�4;|E.��Ѹs��:x�Lk8�e�$�ӝl[D�uJ��P�y*!�2�o���