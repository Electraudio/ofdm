��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�tC*,-�����i�\�}&���q�2/x���b���.+~�8�.�9@��bc�����Q��=�K�&ӕ~d���b}�G���.ֶ�Q��_�e+�G��t��p�Ag����P�b�ý�\z[��A�(T�|!T�M��w���"v�۱NN��U�'Z�µލ��y�[�K�p[&$����?c*-Ѩ����|2�+P�:xY����T�Kx|��Ȉ�T���V��ɀ\�"-&/`��AD��o�И���e��ċ�^���2M�9O6rE �UDc�>]v"n᪐�Ճ�f����C�-�>���7[I/�`�]���DW���P����������}=�a���1R��z�Z{����m����K�:^�{t6��@@RLAƵ��A#�6B�A�xl�vP�sƍ����W}bJ;o�?y�i�G�Z�w�,�|���.��4������Ndg�t�����``
3,w�ǍZ�s�NQ#��|Ԅ�r�Փ�㚻�}v4A�۝xh��a�&�o�z$ ��,V�Ʀ��V��G�	(���́X���exg��I��sO~N�h�]��Å\&���G2 p��5�Ih�[��10��*���g^F�-�>o�^�����6b<�#�����_�J�R��<�����=1F��Y�۷�$��y,C�����̔=C�z"R��^�!`�M;ƅ����s�
���i��+zp���؉j!ް.}<��TIsS��ݎ�����;�y�0�������:%Ť��v�c3o�`"@#4�5��?+���,ھ6%!T�a9�ѽ�9<Gy��}M�U'��]�m( �M�����ѵc�KX&�L�7����y*+R�0�_�աS� >��:��fV�� M�|�=��4�N�i�lI�.��U]�T؏�"��W�Q4K
jl����i����F<@�΁Q j�:�vi�.@�	n6r1R	4����?��t��J�j�.�H+Pޮ�!�z����N@�|#:�T�:�;��tN���2K3J�B���U*�SYk�rc��!�P���������b�G��Y����
.
\,]��úT-H�;u��*<)kH�U[��p�M@�ۼT��0��9��MH2��~�����U�x�p%��$��&����p���	���dj�rp�*)���,W2=X��H�@���#��E3]�տ���q/�9�H�O�1�7Y�"Fك_r�#<О\L:f_+%��_��3�	D���.�����ooX:Cz���`��W #.�wA�җ�<��D,$���QK�c�iT�~t�d��[�t�";��o���q_%+�2n��|��.Ke%��yI��l0TA�����Ե��"㤻����o#`�aPK�Wp����Y�X��##2q/ ��,-���,5�C�7˦B�E�1]��ʬT}J��&�%kT�Ky>��l�W�l�r��\�"!h�x	��@1S�R{z��Wi���i� փMIq+�}%�BkԷ��/&�~��^9�F���=����-�_�?ZyF���@\ޑy�� �iF��x(\<��ir�q���%g��"�����z�r<]t��1e����	(@�+�rQS�p�i�Gfx�Z�j9�� �=�/�R|�J�W�D�^@����ݹ�^T�2�k{�F)��Q]��#����x��:�&��
td,�ČJ�\�~U�����JZ<�Oc���Q�>�v��ɏ����xdOb|OlNU;���+%�%E�0���&F������}���A5�0pL��h\�S}՞rf� ��'ИpED�~P<���w�X[�-�LC2�sN]E�{�RxX}�9�(q\��V��F_eX	F4��|���U����4#�{W%H�,���N ,���*����D�D>��p529���P(̵M��Z���˰ �i���*4c��������ר�y\�T��`�kZ�ub���aL:�#S��<��`������:=��Aֈ���k�����G�����-����r����]XB9�$�dHK�XI.X?��ǒ�tm���j*X���:!��"N"�=���/h\J�f�!���u`�Cq-Z�?��sF����X��Z�Q����z�N֔͝�כ+�cD����@D?�D�1��~9i7:��d��Ij}��r7(0�A�����Q,����X�za"0PMXuy �n���%�B!�`3�`�A�f���-t'��|=��X���)�2����P��D%�Ā�}�΋��@A)�}s�.���	��At�	�Z�6�K�V]�]��U���dx��]����c�X�&��N��ﴉ�!0�^�K�c��P�g[�5�e@�Rߔ��$�=tv�'!wEM�ϐ�F�	I�/ߗ$��ߋ��ϸ��I��}|!&�x���Q���Fz�uk����9̾^�JS���(ulʇ� ��ą~�Д�����+w��A߶�U4�h
n��n�j��5���G��u�W���6&��^�;Ys���\��6����)5���f��e�)��=;�JSm��G��|�~*`��w�)�t�'�s�?��5�0Mx���a<���&�!u����Z���$dȒ&�8��ڟq��mZ�ZZ.��w������T��y��gꁲh�H��?�J�]x����(������sq�P8�hXS%9h�s�up�	��st.����L�i�:�tZ_����ʒ���1�ƽ�i&�Y+��J�I��-7�w�����9����<ˬS!�rv[7�����ݭ*vӮ��y<�a�{�>�-5�����.��MB�_�	�zO��Yը�Ҷ��z2��I�eKG<���ʘ�L�`8*j&�r&]Z��b�>Ê�#�m4�&}��l��5t�0+�8����%�n�����������5��g�TfQ&�-O���VU��(�9B\�D5sc�kǟ`�D�8616�W��Ř��	��(�����o��㟗2�ճ�z�|����M����wН�ٞ@W;�Sx�~�D�Qb�ߓTC�"�����<(�\�����4�\M��G�LP���Z���\���ǌ�&8���;_��<�cr��	[�q��෠N_��,����N�cj���ܞ;�[�ç�D!.ko�D������ȑn�r���o�u̟�+Z��S���(�\��ϺD�a�i��j��񻊑?xܪ��-X5ݹ�����i�1�U_����<�>