��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�	��t�q��Tj�����E�u>�ET�Uj�a:W0�{E9�0#v��g��_e�I���7���eW�t�Z�.1`��u'�8�7p�b��I)�XO���n0����߲����7ɬpÝV�%�T�g@ ��bٺ#@���&պm/X�b��XU�PаgEn��8(�4kT���(F)C�)�@�ޑ�Um-���T�56Xj�}�ڴm�nCO�8���t7ྋ�ߧրkǎ~hc�U�.sТ���?��yk�0���)��I!��I�>��Ўru����}���T�-?�"����$$��%B��/��@� ���}y�ܞ0h㷴�<|����G�֢9���n<��|��X�?k(��x#�b&��ӽ^�,ܴ���X��jNȺx]�^r��`sNC�GVl	x<9L�_4���أ!���m�So#�r��vK|W�S�a��Ѿ�U��<����=�V ��m�r1��&�4n�>{�6���!���֎ϑ$�1pQ�I�'�<��>�N�R?E�U�e�.�\��n
���SI�q5�;���3�?�n��Fh�[*�3�`�pՔ�Ya�e~Ù?1�&�8��; �+��v���zXǡS&�p�wK��.v+E��F�-�g;^@7낄cqif��s��p,�'��L8K�^%Tp~$+4���f�����7��(�� �|6?V�I��w�n�/~�ې���׿I���z�y���h� Su�AШ�ݴ���ٔ�鑇)���K}M"oS'{iV�|�ŭ �i'T��O�͠h���c��#:�!�~>���+��RR�����g�<�A��?�P´3&��T�Oai����ND�Kv6����
f1b��m���01�ٻ&�6��'݈.B`
�q<<��Q�$i�������z���Z�K?v��?6����}�1�K�&�xj���z��-��Kn��ˤ	ڢD=z�xIc9}-�wG#��?�3�|z]��To&!��n�����6�/�{��ކ*� �m@܋��J�$����N���%g#��18ƹ����"N���~���l������Evd�!�g®���WL��H�R�`+`Tc��@�l�۵2�cSE^C8����-�U����&�|���|���{iC~�dy��_(�({��yDuy(���aqY�D�!����G�C��w�1>Uoا���ͨ��_�/��#�{�Z?Ϫ��]T�(r cz�i,/#|�_Gia����ŵ�D���ia�ӫP����^G?b��j!�����@r���{���/{Q0�APUn�C6��r�j����B%ar�M�u�!�D���u,�PCm���/M�I��z�ؖ��\7{̉x�Q�B{@��}�N������'�K�+9ES@9H=Ф�J5Dd��U�����3������� ЁFˈL�q�,����jR�k�pebhnD(���1$��V	Z7*D�D��v?�I��� ��5���<��_*��G8b��W\K�@+�����hK�;j��2(��ZQ����I0���+X0N��D7��)��Iu6�5y�<o��`�n�s���4⻥�
Y(��v����"}��'!�F�vB!Hx�d	;|c��}��;��ޖ��t���JMM����_�+J.�_�z�z�f�^��Q���D����"�TS;� ��};��Y���j�P-#'�9��bbV�R��'C���|Q#妽�r؍�!�ں��TL,�2D�ǡ|H�O�&�!���������V�P�-���bq��M�/�	������l�٘[=~Y>���:�I����+�nK�="}��`�Ί�4�T�|�L�5�H���DY:�z�r���(�4`���`�sl7:G�u���k}���c�ɮj���n�{�ӻ��Ϗ����li�b�6<G�*[�mꆭ����V�z���rP�<�}���f��\��Ӫ+@kh����0]^G�
�Y�b^���:jZ�^-�f��Q��;�zg����n|	zN��f�D��.]3F"5*�Ո,�X��Up�������VŋZ�����5���WGs0�%�a#��<S�H�H�[7$l+��r�� ME��r�/j.�・�1[�ųI��5(+�Ee��/Q�h�m��CXg���[W�� ��/X�/�,p#S�W�ͨ���Z���Z�(�/��|g�9�6��c���2�����!\�ĭ���Κ���6��k��G;�rg>��M]K[f�#�!����iA�/��=�THj��G|� ����dJ%�uL#x��%�E�i���U�ԣP��{���#�I�Z2�L= l����aj�����΍@r��ԏ�`d��5�Q���4��ǖ��Gqr�p�s�W:㖐��Q�u�:��&��=�6����N��8<��T��	�������"�g�߯m��2�T�n��x�*�A(������>_ ��Y	��D"�a��H�Bʋ�C�G��&����9j�;~�0�E転���B?�\o�N �2�Y�턮��UP��+g��#;���b&{��T*����m(}�U�\D�x���<�c1�'�
:Ҽ�9͵���6��X�����^^���F�{�{!iZJ~����i�Nf:�N�U@($�!J�:uR�;�z�(�\���q`�ڧf�DS��nXŮ�G��Ju�8�`6���K�+�u�6Ƣ��Q���SGn�#s��* �]io)�Ea��}$��PZ�8e���hp���z�M9�g���^���w�P�ܙx@���%1��׶�L�X����p"F���d�a�d�B÷��ֻ�`/���:�1)ą��@9��@��(�5�
��̮�D���N*��^��A��b79 4xɾ����?@�2����/ �����֡}x~�t��<��V�v��1�S̳��ڑ]�U�lq���X�Ȓ�{@�^k�ڟ4���#�)�w������ԎIDf<��,L%A���x�r�NG���m�mFҚ�_.��@9�����
���@S�T{Ӿ{6h�I��i9�ҧpJ<U��5�u�Ҝ;�].b�.��ԍ]�&P%��zhA��Q�x_�����jV�<�gg
�"7�)b�]G.�	~9���/���_l�ZL*�2;��QX��~dq.E9�B���Jj&�PW�La
8�����%�Z���f�o��&"�i��1 j�1�N�!4�� ��H�����Y��2����	��(�q��%�#RMã3���J�9�g����
D�P,�ծ��К��=��u�(�ӆ+��&����Rs�G�4���Ut��2�p3}{���20��6��3�F�cku��;h{��`Tv��]���	���7*�f��Q���c����]��]E0��~����L��x�jp-���in�ǜ3G������m)?s)��Lbf�e��Rycz�CĄ�����O��ʨ��Љ'��x;6ba^�p�o��V��m2�D*[#�o.+��E��޴v�b+T����ֵ[A�����ġ��`Ϲ�>���u�El(�R���CW�0C��~}�8,��yv#@0e�L��>AN�09���1G�2���ŝ�]�8��$R������� A��$�-��̬�_����z/q��p�E��Y�⩣~��N���*�}S��j�BmkIp����83/A>9IqU�A�l��J�#�*h���r�N��st��x�&��1Y���ҴK��[;]�� m.S�T�y���{l���BEZ1� �0�9!��9)�~�5��`ڣwt`��/3!�lP�KjNb�h	@�O�u����?L��s-�0�1�(>F�S)U,!-Q���9�yb�BI�Y��̓��q�����|�C2�Ϊ�U��Li9���n\ I3�ƐxG���;��s�n�h�q�+X?>	~�C3U��X(�qu��t�'��k����X���ճ�}=�2Xxo2��y�N���b��O���P��P\Y4����p�$�M5py(�/b�D#d`�F�r��	�ju�|e��A��bz
���,1m>g#)N_`!z/=�s޺��t�VJO����aO��Zi:h��|��\���{�e!�96��dl��_�~f �ʮ�Gَa�pV��SUJ�,˟d���\��ix�K�_�����Ch����7D�,�H>�y��l�-�#�����W�ݶ�8
���e*�qAե��@�̩�6�]�s5����*�k7�EE�v�K����KO�2���I��7�L���Rq�ҡ'��c���d��<F
+R���{�/��=<_�`��a�Q���J���Cq�U�9ҕ�l����&��q�� C}�.S������t�#.U���Y��lt`�	�� �����W/N�{�_*���wē�$�|
(mn��{�Bn��1��:4`�V$	�6��q�U�nO���/׾^��}<�sEt�eh�`��w~ځw��TY��{(r���K���N�5�W�����dӮ��t=�E���VPp�躍�=rzJ�;��Y��	�.*a�RG_��a�tD���d��Hz�����7!O��R�t�T��7|����F��L��x�� �h��I�ʼ#�@[�%��K�O^���N�Qqx5(�K�F�%��x����mf|�J�"�y���;��l���Q� �+)���Λ=Ʉd�CD�\���(�}(d��5�ׅ̔A�T�'t �ߋĵ��c��j�ټ�����[�{�(�'Z�1ƝC(5��o�A�.?�b�E%#�"]vxzI1/�&��V����"V�j��b��ۼV._w�S�$ ���ž��t�g��ܪUy��F��	�b��٥Wl;+;�JbԈܝ�<�E�\��m_Fx/->h�b�UJ@�ж�.��5�%`��3
:���83�v��I�(<wxWܺ����]{ j�?S�Cq`��� D.��I�dg�2y؛�@�74�z۱[���b��ެ�o۫nɻj%8'X�fe+)�q�R�����yה��,qE�8h��D��2nt�<��t����,�� a4���<Ǩ;4@ �hv$0�B��\u�@�����DQf��CgQbզ�2���r�v��E��&��O��A�X�җU��Z<!iV9�m�t]X᭝�|�䪫3np�I���E.�z�l[sE]��Fh�N>n�28�g�ܷ���Ƽ%4xn��Kj��(�؇�h�n�q;
iT�7�oq�u
3|�h���ץ
��qa����70����b�q�"�0�L��"?d"~��^ۓT������=jP�1P�@ 7�Ň~�ڟ������C����p#/e�������5(N
,.h�Й%��8"J�Eg�ӧ�u�T@!�P�!.�l�����vS�]�g|�^/DN͖q]�G��s:�S��VCr;v�p<�ר s�Z;!��/��f����~��1N�S/m��#���Iv��9��M��}v�W&�Ln>,һ(�^Qt�
o��(�	kü-���,�${�+���i�V��Ebr����;2�e����#D��w>Wp��Bԁ`��S��}������@NA_'r��\�60u N�&��Y�M���5�2���"���^���u��I�2ӂ�}���<�v:�I��(�PԜ�RQ�`�8~[��0�	�|jهW��l��Cq�7��oL��+��ђ�n�b+p�v ��R�u�UI���)�s�$,��H�R��J�s؜W�!��R���doO�(��o�*�~p�qZ相e)6s�(Po����b����?�l]f�w�;��!4A��4R���y͡}T�`zm4c��Hk�LМ,�D!291��b+�i岝�-�6�|\��K���w-���&�d#c������� �+��/{��"��Nv-xj6N2A�b6��.��������j�c��3�c���o��b�Y�=KOHd���x1=�hYT ��;]�h(�l�<E�,��c��"i�B�.#?�D��Ը��L0Ԗ�H�"���+��Q�h)j���~	�*��o] �v�Y��חpcT�cvIὌ�|4rq5���$�3��X��!�j�o�A�w��W�ɸ�1�7���<[��� &,6r|7�j��D�M:3&��J�`���H ��~�?&-�86IFݯ|&����؎���C��:�S�K%��=�B�K�!�x�lu,��V����������}���NG���
GX��2fP����9��o�*C���=r?a�0�������I���ǫ�� �uX�,6�u��V7��f��,*m=��MW�!�2� ����GDϫ�����0����d$U�����[�_n��b�F��Q��e2_O�GQ���9Տ��������i���O�1��ޔa.�̸oS���@0�'��$�ige��M���s**����L�&Ѕ�jc���D�@�����@��j_�AU���+�c�m8���3�%��p_�f�`̷.��
�#��Tq�q�����is~�[��o�e��1�1�ͥ�`&3�����7x�ވ��.���.|W�
c���֋z��Z��k
P
Ȅ_-#ț�G'	��{l�����0���1��Њ���!,؉^���e�@����,�/W�vT�A�0*H^J���J���R�M��6����=3y��Y��>eB�3.��j���l��/(V�S��k�	� 8[A�Pm�̝ؿG��s��Xz«�p���t�mKSүM u�Ž]󭌿�?'�&D�i������	P|��l����V;�FR�O���@���m�&�Q�P�m'�|���ti'R�N����
���ރ�W>���a��öЍ����B#
G���Zp)4:rC�uCt�����R8 ���4�3�����t���rҁ��%�
|�6-nf��4�Ei�P矋=ӰiJ��u�UD���� 9���42��Q����(�+,�t�z��{,NG�ȌY��aJ�b�"��P�`�aQc�ؖΧ��ϯ�x��P�\�8P�f��=�Ɲ�dB�{��:0[���	�43�a�����;�2��3���`JVީ�l�F@���l�7bc�!y���&*8�^y��D�!.\��o�l����_e�� :�| U������x�D�agG��a2�]8z]m��'w< �A�1�e�W�
����ַ��qY�;�Xڳ�}y<�����Q�(�:�"��Tn��]���Δ�A싇�@F��753Wo�O��X��b"L��