��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0�+(g�>.b�p��Z��N��]_.�c4�1m��}vKv�ں�ى����LY����M�ﱐ	ٳ���08֌��@�G�Ȳ�fW.���9�=l99�%��{�J�F����L' ���E���x�g���{�T��;]�&��ӭg��Ӄw@��3C]$Ō?�>��
�m��pr�����[��-��|m�zs�!#����tZ$w�»EC㇥`%�*�V�W23C$Njp8�A3珅��)~�� ?x���>�vL�M#n��w���A-��7��vg&�da�+�(|$�9���YEQ�.�c~��n��5�T�z"������p�3xsɱҤdUj���]��d�CXa��Y$���͵Ը,�%M����o����3�l,��L��Ur�MbNH��F��b��ڳi�W�zy���уg�X0�*�(�*�wC�4��fO=v�d����[�
��;��RR(�f~�~���A��IcϷM�7�'�s-�X��U��4�b����]�-�
k��	�
��bv����/l�����Ha��dM(��{;ET�:�9�;7��������"�X!b�m�y�&��S���@���� R�(�Y�ʜ��(���|ǄqE�]1V��R2��3�����;c?��V���j��[r���\0�;,���%T��oi:�
]V��޶�ԛ�ƪ[�&S�S�[zX�W�9�42x��8~���^�m9�_:�n��#[���4�䧩X��onz7�X�>�H�9i���+��'* �*�}�It�^�Vg!.�}�� b��(e�3WR������bZ�:���^��|��*T�q�����Cu�]kĐ����_�f]�ݬ��i�9�8������ ��Km ��D��-_*o����&�VRV�VsO�������Q3�O�$�Z��餩U��XuX#��+�>�?�� ���m���(���$HPr�<� �������Ì���>d��0@�$�:�l�;y(ݮ�{���}ī�$h��_92(�i�Vs��t,�3�E������q��ſ�yh�t�&g�$[<��j)�����\z�nC����s�+[x��͙�Vp�=��#��F���/�=C�U���[��7�Șz[H�
ɳ�c�9<_�lXۛǹ��v��%�[�a�c�)�c�J>��%LA��ϫ�O�˨�i,dT`�G-0Ooo�:���i.fz�Q��s�}�7T;�Jmc,RcD�o�a��
�-n��T�R�j���T��qˋ�M�Jk����������dX�匵*Bcn���Y�G@����Ӂ� M	}�}���ʐ�[Q��W�-�Ry*�7u��C��>g�sY+��˶�m�fvF�8Qvj��'P~�,�nw�F�MPA�����x���i�M7�:�z*�����t(�Ewy�:-�yLF~��+��Ror�+2���l�N�|��XM�MG���q�Z��6'�����5����S��+��u�������R�ʂ������z�0��=�[��īm�����p�}�8ܕZ�"�e�g�>x�Xf���z�1�[����#�seF�{ܠm>����Z�TG|G¬�~�>��pk���Hs 孎i,B����>4s���eH1�ςP�Kb�nc�n��/
ų���+U5{z�%�I������_�(3�ro_e�j��]���l�j;���"z�����N��Vf��$�,�LSE�HH�*�t�����j�:%!]'ԙ���0
�k���{x� �°��4�G���|�&E����R��XؒV΍M��b�p��@�:4�T7�S��v��-F����E���쑍����c�J ���X�?��}�'h�\Z�9�h�����]�!�18��c��㻏�Y}GKU�?.���9��E����z��X�7�Yf7i�E��D�kk�޹�&}	�%uZT�� �yc���X�>��ġn�I�"����Zt�l%*H~��歇��&�+���n[��T�W8��2���1�#�XC5-A��9T���y$ܬ�,�$�{XRҕΪt)�Z�>�����������y߶`�,\�<��*o�{�fty��O
��w&-{v�m\+�z֟�j1�%�4���JM���>���bƠ4���c#Õ�L G�D����nY�N�����R�ܧ��6���Y��-�U�T���N�/[Q���+�m�6����\Eu�D����]�M�I�!G��/�]+i���K@k�����O�oL+���aM������I��W��_Q-t�f��������c~s[����-m�L�1-��6gH<Ə�Դ�6�& ?V�%��TR���M��$'�;b|8�!�C�{�]X������c4�F�n��W�'U��NNbL!:�%t��3O��?1���ٰ��ư����O+H�����IP��p�F��??���5��],&��f�Co! [���~�[mfk!��a�c�I���U6RN�*s)��:����G;F�DpT�¦�|?ػ�i-�=6� �I!����o]������[�ӜR�Z@�0�l���K�Q�2p9�%/\/�����7#����_��08�}4���Y6!�x�K�x`���oD{�a�|��#-x�̀rK�R�
Z
`�bʑNr�]�S���/�M����f.!�ԞC;u��YGH&��s�ZT��!₦�렮�T��
%Ma!��;}*ൕ\����i�w��}�ޏK��d���h-���XF��V���;c'�R�����`������o8؄���:����/{eF^�_��4��[T`�Ї�:��.	3ZE(�P�Mn�Wԟ�	9د��C���)n�7G�`DpÊ�C��_е2��Z�b��!&�7?���F3�c�1��&2�/(�U��қvH�X�Q>�rߟC{�X�GX'����Qd�<o♐=���-Y�wcGhd��8(YX��Jo֠ŷ�
ҷ�f;F�l���'fޝX��Q��������S���?�D�`!�W�
w�!S�g|��Y�BX��{w 6��+�QhC���h�i�L�$��@��w�s��Vj{�q]�������&�8�߇��)x ���;I���#xJ�C'C�F��x�8߃�s�}kH�>���h�U�쬬T�5D]Z�6�;��ڰ��<� *��������hn�(�g�ֲ � 2F%�1��fF�L������i�<}���>�^�e���)$��v�R�P9���]QA��뇟�`T���(.f_�O�glu�DÅU�����fşm�&r%�a;7�ً��D��6��]]1�=�҅#�])j63��0H��)\GĔ��.	���+l��
�Na8j�6�r���M�8ΐ�I�,�j�R�[�'�g/�}g;E����N�r��>�|`��²�e�0��c�BjBL���Pv��r����/�o��73ލH�)Ä7�y��6l��J�Ɔ�����\�K?6ֹ&� ��!ڜ��v�pq�O]`>C�B�|�<C Acf�4�*\6p���+2����Y�	�j��1�ɷ'� K�8]yK(�
�e��9�����[�s���H��`�i5aL�����u#�o�>�'̓�'%l&������stf�8Ҁ�����B�΅X]o��Y�������N�f!�@^��	�ѱB�.��ʛH��2�?�%�=��}�������r\��d�_ci G�Ӕ>�8|PsSQ�9-W󫬎���qlMo���f5#�Ω /��ưG8�\���
�Ó��>��!�ڶ7W�M�O�l�%�KnǊkO��_�Gw�X��9�Q��)G�睸���5�+p���vYȏ��Y\��H��9vyg7~�PV�ex�Q6�Y��u���Ĳ�Q{��_�*��+*��| �r�0i��^�v���L����=�F~UW�^f��:ӽu�O�w;Z����B������b���or����U��Nx�"�B^�i��Q��8d0��o�k��f� ���B۪�Tܜ�E�bt3'����y��Xh؉2��VD�u6�{������^j���Ȱ��	����|�X�y�}R���j;\P.�ǒ�v�J!��)^�k:�U��.Oe�O�PYK�U/��<��*^�;W�i���m�3"퉾��[*U�F�}e��Jr�r��ٞ�5U�������N����}f�H��Y��3�:G+��gC4B�k��C�*U�#I3���-ƻk�6�|`d����[	`W]�a>dQ��Ϟb�)�+"��_D%ۑ�*bLt���?�,�č�? =�����J��J�t�x=�-X�5Z�̝�����qb��Т�NK �GXc�T���[�@b�I	�x��(���/!�_�����Ч@c���S˸�-��2Uθ�r>�vB��889q�.I0�����
����գR��\cY�u�3Mɞn�ِ����b~ּ@�?J�Eݾl��*�g���'1D������R������LI<�/W��� ;1��@[x���#��G��y�f���_�����;@)��L�ނ��Z6��1�r�3׌#6_Ã��]�&�L����F���H��Ƶ�*�C;b]s/�U������Q���%U����%�Q[���D�w�i��Y���z�pcng�#��[v�?`�	U�@�����\�����h�����w�����3����Q����X+WE�����?F �D�]qB����L��ZFo�Ws]\ >-�%�l��֣��z�I��a�6�f�����8?ܢ�-��������/C�ݕݙW�Y���xߕ5�7��	����q�c����� ��%	�'�&�ɠj�M������Z��'KܔS9&��V��z4����4�{��1-x	�&	b�f��yI��,�4R"�T�ڊ�Kq���_Ƈ��t�扉��0����t�WS���<�ń$�ˠ�ޥ[��K޻��㷃{�L�Na�!�B�#�F}Lᓚ6Fyy?#�0��x�~mV?�'�����i�v����g*�|��ur*t)�f��E�[<�L/�
�h��b��k�1�憭=�(E�����"<td � �[jarg��DBz�5d�5�n�H�9a�ǊOY�Q��9B��K��T��ǈ�Z"�;{���h�N�Yƍf�r*�\�K���3�m��� �@<h�#O+9$�8,}LD��q�)�C@2���p������H�l�a�&��+���<�W�d+���z�蹈$�G"�2�tHB���������No`�+���5e5��0��|4J��_;��c۲!a0�\�)u��0�Xco�V���6W��e���K�g#Om�A�lр�;H�蜅TU�"�XM��WWW�!�}!��܂�5+�=15t���U�JW��F���?�P�`Z�(1j�Y�d�]M��Ԝ>/tk�j�K���Ae$���L<A��}$�W�2΁=&X�\mP-�g��2 �(δ��\sR�ys=�:|�6����ӓ#�o�� ��׼�כ��h�\������vb���L������k�����}�'}�w�r��-�`U�ȟ@櫫zHdu�f� 	d�0���k"3��B��I�m@�ɰ>�N��.��P�)~���tÎ��z�j2M��f��ϊި��$Ou��u]C��g�pR)�_A�F�[�������o�q�[����X��J��,�����Oed�"0>;�v�қ�D�m�Qٚ���ՁB��%Y&ݔ�p�
�Ԍo	��(�3qr(�ˊQgɦ����T��f�iw����(�lD�W�<g����E�	1f�� X���t�%�!g���	��5P����F�v� �6�QZ�']�vK`�
�6��%1Ն1'
�ˣo>�e��*hX��E)Զ f����p��0"ʭ�?~��`���]��>�p��K�\�c{�0%�����-��o߀Ŧ~`5�����eG�W�ʹ�������'g���Հ�3g4!��(N<�~��&�":B+`[��e�0խd���08|��hw��֔���m��ft��P�Cc�{�r��>��T5�Eqg�#��ZK�����%V�Y� NwMZ�>9��v8@�z�&�Pר{�Y���CS�������X	��G���d]V�Ǡ)�Q嗻2!���M�D��ź��	_Y��)���6���Ƚe���fz�$��0X�Bj�˾�����=:�ή��sL�A�V