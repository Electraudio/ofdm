��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ���9Y:q����&��q�h�-������AwrQ��R~]]D��<��+�<d% Ru�'�X�?1��T�"�Isz=����$��n��m�=�����*��{ _-I�LF(W��&t$�F�eAd�D�P��B�0X��#�Y�z���x��y���ͣ(����(J���ߜ儣�I�ݛ#�H	�V""�JC�,f.�ۀe
5�}���7� ��x�M��i2y���b��Jڳ?V��J�}x�Cr����&�;�� -n����>Ўy�>]��(�S���̬Yh�{���;��6K1�Ÿ~�0��0i��K�s�C��g`��38#�f�E`�5�����%�Z|$�U�}�V�U^���C%�pȺjN@ĝ��3U
j"�d�?WcR�I5i(W̍��3�d��ǯ�5�9~��f�[���S-��u��>���h!�&#��-����Z�R?.�r�f�[���yW��S����J��=��z�L��C�gXG�����]u���o���]�J�
����<HM$�_��p���<�p�U	�w��T\�b@��d�ʡ6mtz�%�U
'=y\ �x잶bGWl�K>�xmM�L�nRG?�;��P+ �����K%9�0�D�ʭsf`�`�z_�����I�T�v��٫q6�(Rbۃ�央T$�ܢb4���o)����tq��;:��8�
䭃����ƺ\SHŕ��$�2��O��F�x�8`�E�^�N.��SD��unI2W��:nKf|��x�����YM����ó|�`|���X���]��ؓ-o��=�[@\��*��_��c�����Fs���/��V�~oCl�z(���[څ��l�fc(sK�@�����g#q����x����?�C>���X*�Ѝ�e]�������3���\�E����r��fE����S��ҧ�~!�˦y�':��e����#a4�N�WPҠ6�x�Ju��`��g�ɨ"#<[�k4_w��y��2��ǭ�,�us<�E~�Z�(�b`��4���"H��S�x�uڹ�B������=�꣍x�cuF��OZ���Fpb(#�����x@�$ߛ%��8��hP�g���b��펴+��V���Oy��[ܦ�
Y���\.�;�ķ��P��hu��5N<7-�?f?�R���o�6�>��v-?G/�x�s��a(BŃ�ڼE��X�$��x���V8�BXZ�R�P#�.������Wv�xH��8�h�y��K�o�A�t�xFY��"�N��h���&|�EC]k���?��"���Vd3��{��߸��L*p�^��0PA���{�C�Yh�We�x�K�d`U�|@��^���2D?��ļ$��=�.0���EȂ��ު�	���1}�W�gݲ}8�~���ǒo�*R�{��rd1��r�8q+�pq� ў�����}̳��F�!��c?����h�ʠ3����{8��z!�w7��*�v��S�WV���评���F��Ɗ���$�#l�����������j�:��!�F#���;��h<�\D��iz�[�"�'�hoൗ����T�[�n"�S�sѯ��w��E�� 'Fi��1�ѣ�*Hb����p�r�hгUX�7��-���t䘗��Y*F�8ݰ{�|��L�歲����Y,��s	�����Hp��AH�W�Ϙ���=V���)�U=�����7��|O=��:�D�ʘ�Q�Uܞ{��u�L�Z�O��:�P$��f�[��������gg+tQ/-@��c#A�
�F7�W�\Z&F5K�����/�=��<%2��g����)���CÀF�%��B���.�E�]se��a<�gl�[X,s!.E��M>ڡ��Ӫ�2��Tw��Hs;���[5�◸>_͕������ȯk,KV$������+��R�\<��}P	$l�Q��1%h,F�Үi�����hx������m��!��ި:���!t����M�*�᳻'bT�7��)�ҝ�96�4��6�?���/N���2�,�� )bj�}Y&q��i(�y��.{�}��v�ܑ�%3�n��k�O�e����W����<I�G9ܒ���.��c�����/��3���#�Y��B���dv?��4ӹ�BY�⸎-�>������x��ʥޯ���� ��j�O��0�TڛZ�=׿_U����eK�}c��`ч���~<$p��Ch]_>�+�2d�xר`4����»ʾ�[�Y�Vy�� ��2(��Ǽ�=�s�v��+�����m^�^3tO/ȉ�oo��uG׆Ay������h)�|!�B�AQe�ܱ>��rd���n2a�[�s���dUPSgdy�I�gĻ��� Sx#�L�7�1D%k��:�N�dH��>����l�9�7o�`�ń�i�n��[�m{�x���Ș�0�ҽ��ѷ�*.tEv{(�����d�S��O��Xى��3&��ng�������NWf��+;s㡣�|��a�X��ְ�Z�����̋EVct�1�ZfȊI%^a|�	�P,�I!/��}Dr�]/�6_J��^���?'�?�}����IM��c\f_>'�p`K��k�Z斘j $:c>��>����	
�<�I��Qp����{��F�}���m����0��dxK��>2z�K?���Zw�P�KG�cD$�4��J���&�?46w��:,ې� ���Q΍J�IRXA��iK8���d�oT`lAq�ø̳��� �G]k�׿�9P4��Z���>����l��'Na��Bt�\ڃw.oLd$�ms&XZ��.�y�H�S|�2�gӊ���Zu���3^+�'ޭ%���/P���t�ݏ�H��zn�����go�ȱ��B_���<bd��RIF2K���$]�� g���U9��k}���f�D;`�C)$F���6�.����=_�iω
�"�m�e���q7��R�7�g�Cza$Y	�Bj���x�Ѽ��݆�7���E�n�~�-S=�����l<�o�)�.}yE�
H��WQ�⓯�Ֆi����5�]�0#p�o�)�ݣ������A	��<���9�b�C[��&���Ѡ���'z�����n��\�pn�{h�ˡ$q3���_f= ��H���fy(�r�T���N�m���lI�	ᆴ�;ylF��� �R�|q(���J&t�Gn\K����$���8�jbB_;�/Q�n�\���΍�U[K��5�[y�QHW�f�.��������+S9iv�x*�c���l6�ʈ�p���QӦA��3z��k��Q\����AI8����q��!͚E��̘��6Z����['�{b�����bB�H�G�������J2|M$6N�u�k 8vi���+5��W��ك����A��%�vO���/BA�+�jj�a �X%d�'�wزv�'�j�ǫ�O�p��̗ Z��ɟ]|n��� �C?wP25�G5ed�?����B�Z�g2�8\֟��	��| Pf8�GM�HXpP∗���|�&���NH��Y}O�W��z��������k4�d��E^|Q�k�Q�k������%��c6�֯��I�іY����\�eaB&S6����V>��l��t+��S/�ٱ�����J��,;uZV��!r̶���5��i"�wմ��]������\͍�V�TbsM�t�Ez�~�5��Jw D��vC�?x�R�ۮ�:�DB���q�w�󛵡R\%��i�X�3��8AM��ge�-��ӂW6����:{ ����A��M}z0�3=�g�	��Ż���&�ސ��#zI�.�;�Ha?�C%;�Ιt����,D����im{h�I<h,߬�[�����d���K��W�=�$.#Z��E�G� ����S�O���DHP��>����D�8�=�6x�5UJ.�'L1"1�W~UEC��m��;l����LP.����J��Q[O�Ğ?���Qb�^�ы(�od�+����n���@�u5_��L�me���{���9Y�G1�7y���s��:����7�V�gv�;�Kh Hg��Z|�'�V!L����l&�%��1h��V��0Q���u��oݐ�,���Ҥ¢��$������D`ֳ<�����6>)�vio�4�b�.��V�T�3���(�+^�x�d�G{�ʝ���!����uhT�S�)	Lu/i�Y�o[�hXPJ��l]�)?v�r8���9z�U�&��4+��Uiq&�"&�7��V��yJضߎ�ʁ����mP��:x��@H�G*���'~1�-,9wY
T��H�iY\=M �}҇
C�f��2�p�- BT\��RR���j# �;Ue%��-?����oY�6Y�׾��s���Կ2G��s��������޷~��`"f���M�qX���'HI�VE��h�Tr�CÃ(�����zeJNS=}5�O�/�!=uKZdk�u l���ڐ�6�����*)��鮅r�g�Q7Us�T1����Ӡ_J�]��i�Am��6Tč�oU�co��xhS�-�*.n��_\����W����Jkw�| ��<b�69r�5��ȟ��_X_�@�q�J+��.�S��aߋ�s�\y�B9 ���9}�s�����U�-	XߨiFA�X��}��
9����-X�	�����@6����P���y��,�dl50o�!�N9�Vr�z<Q���qm@4���%���+R��;%��gXk~�$���䲝t���H�,2����JyZa��F7:%��4q3p��P76G}��9�h*o��k�{��z��H4�ر�o���;F�x{%띨��&ڇb�s�=�Qb�_d֓m�<�����3T�3�>lmm�}�}׌Yd&VNBi���|4�b��T2*@nT;�JB}�;���:�s��Mj��bb���:�ԛ�����Q��C�w��n�Ŵ�]��A��C��1)�'���j���r(�����a��e%P�ҁ���/3f&mp��[���7~H��\Vu0��-ENLZ�[s]������k����ٚ6�9��0�V�خ0��&G���z��2�KװV�I���<:��@o��B� ܋w�X���#�^LH��m�W�X��e�ͩY0;,\�P���!h�ڗ����^
=��X���y5�%�S�F�1k�C��b�����[�9���<8�IY~Ӡᐼ4���J%sG!�+EԚ�o�$�B̌De]"��}����/w�k���.XG��]Y})��ז�������.��Y�ϖ`m7����ױ��:vzTl����dq���5�]�k�M]l��b!�x�?rF�	�{7���^`��.#d��f�� {�a���$T_�E��«~�	] �^�����x�ESe����/�U'���5��S�p�G�1I��.��k{K���E��c{�ޗF�㿒^32ĒMcű�d��+<�Ð-g��d-'KM�zX�W�p�5��h'�/]^x�\��]�*�;���f��6�.���$tE�؄�a/ʐ����b�ƎMS��"s"�y
ZV�&�A�N���!�� �2�'3��-�[O|헄�Dv�(��)��6���y֠/G�.?W
��e��4�k7d��D"�S�$�ι�Q�B��H7��2�)�e>>)����ơ�dD(.c�,q�!&����R�?`�8ȁ�9����
S��C�#/��^��.�CL)G:b�j�o��\��=�_�ή���7s<��X���I������^���`�\��P����N?l5xm�'f��Ie���J=�=�Q�`����,��Q�>�=& ����s|�����H�;u�(��W^%�^vI������+�;�*~W��0�e��/�%e�bP��7��.�i_6 Ki��b]����v���EL�P�ґ�Z�z�ä��:����]�K��(�`�r�u(��uGq���B�s���z���C�-��6O2\b9fmJ�˩�-�_��ׄ8<`���+�')v�Xz�J	Ν��U��d|�ԏJJ2���y�̏F�J�uet�C��[����������
վ��&v�.�����n�B�՜��"Y�rqeD}���{5AL��Г���q���x��h]�`�^3((�#,E҅�v\u20h6>�[��� 3\?s Ƒ.C�wzT�R(�rSO�T�>��Lɧ�;��=B-��qr�	f+o�#��c�끾O��,*��Q2�)�8TmP���ݯ����E�Ú}(no���պe�z�X"7��Fl��Iý.$~q.`��r�M���F�z������F"c�T�K(�f!$�TI�����$D�Z�=�i,����dq�������IY�x�ڽ���-H��b��H��ܶa�3$d�#Ŷ�9+M��7w���T�:����쬳O�o;'��X����"Q�\���߫$ ��jWZ��{w=re՟x>�ӳA�W>Ӻ���G�x�~��������/��-�)�ʣ;��d`��
��o]�9�N�ʊ�2��.�;Ew��Π,�_/"�L��>�O1�脸�=���Tt��/QA:F]�þ5��<�޻��y�����l}#\���EQ�դ�-���1�r0��?�L/��;q ~���o&��b�0�5Eo���7�$���&g6qy˦��K>��P�rs�=5��P8����`��=(P.����!���4�>-2��h�OlF@�-���ROc�&����R4P���7c�i���3���OoL�
F�S�cu'/SV��ea����Dϲ���������1�)�8\�9��t�d��)ݎ7 ���]�y˰pQo���2l���X �*B�c�a��%� /�� Ȍ�C�C`�{���k�&Z�P�0h�h��5.�PDOe�?��F�P���p^������"��5"\HL�$������@�87ΙV�㸌��P=����[~��'�0D0*Zf�C��ƾF~�.R�����,���@e�b��r���S	�&x0�r�#i���_�v���R��������.K~�Z2g棵c���dol����5I�����i��GX�l���?�ð�z�ib���n�8� K�.[���[���4�b�5�S=��n�8�G2�Ka7#C�V_��PL 2���Na��AX;I_߂+��𗦢0���7�o�����zQ�z�v����
�	�C)��G�
��5�SW	�ʫ��aW48��޲μ�]����S�;x>�F8��3!���E�u�A�ٹ�~�Ai�B�(w��x�X�2��noc7��W�y�y��P��Y��m5W��׌��d�����~�t$���WlG���櫾����4���L�Lup�%!*��":y�C�|ȡ�X�Y���y^-O^%�L-�M)���5h�hԾ*�s��|W���u�������X��J�}��ޝ�X��\��,�7����0*/ ��ڌ8��}�e�Q_p�����5��+qu<�#ܟ��%,^��0�K�p�xЂ 	]��̠�+l�&{@�m�t^��p~ږ��v1fHɱ�#�=�z���{aR}5�Iin�Q��RE�a�d�e�pHb0q��{���)��Ů�@�a��5P<���h`�p������d9���#���x�&�5�'�3�|��Yvx�BQU��\ڨy�=���JK�h�� &p�V�9�\�k�3Y(m$��$�ߦ?���SXT|�ߵDlYq唡1�D�4��$���0J]Y��_l�e��=���נJ�f�{��%��+�.-��Ұz��p����Q́�ā�=�����V�_��7���M%&ʙ'='��%�Q�+�\ Nv`t�E�Qu�<+A�9yӇ¡j�Hi�|�@�6W�t���!&�z^V�
�=cV$�y��{�,.�0A��C-�=k)��t��f6ì_�[�q��-�1њ�AD����G*�)P�ʷ�kewg넼�to�te?"��Ig{N��N������V�t�8���@�ˀ6DTD�q �zq��0vO�ʋ$s��4�&���_�=�
^l�TF�\6:;
��%��I���ـ�Eƫ�6����`ic܆�+Ol=�:�A�hB�6��C�O�z���Dw\t���J�3~��[���vh���ҖQZ&�b�J["�S��&����B�,wҽE����Է���z<߶��+���&C�:'=�R��<�Q�h˯u��,���֖��/�9\��}�9�Ի�E���[��2�ƨl}��\�~�Y{�g.����� Ē��8��Hҕ�b\���M֧2F�',3�z�7���x�ʞ��Εﻩb,/s��Ob��f�	��<�Cx����Sه�'�/��았����r��*:��/ļ�T�͔�����_iƓ�a�@� u	z��J@����ڀ�]�AŎ�{��x���fp	���R�k��ˊ�����J����^�ޘ�d 2 	�j�&�Q0�}q�-��:�(/��}8���
��[W�E���A֏3� ���<�PUM�O��
��%��z�xH�Ʉږk�.+�.�ޓ�tj3o��D�P�Ӟ�giK�����7K������>�I"ƿX�:1ɴpX�[�4�z�������ܝwvivZ��7eƶ�Ĩ��M������˳��ds�+�u��=;۪Tx��C'h��WQ�G��;B��Ð�ƒ�=��-Ai��1�-�w��F:�QP~f&R��B���\��dׅZ�L��X���|���~�Dl���WU���,v����~��u~�B\R�������L�nOP\�(��M`����y�ꃰX���Z�o;JU�~(s���@z�Zp����Jdhn_�������d�Q�ˊ�Z\��c�̤]
��IC�1� �\��M��������t�P�=̷f\5kV7�-�՘z}�*�Ț�*�9��/�r|�
�1v��_��($7R�rO��T�N^v����x�ƒᛝ�C��� �t�!`||�
N�Ĳ��g;!9�9�r�n�{���z����׼J%�����Gjou
*QE�c�H�{�T�$���/-��N,�(�pL�ܽH�'� Ǧ�9���:*�v��Œv?�&c`F�ПE�@���q��`�l�=�d���5	r_tf�bP/��TOH�U#�N���w��o�K�'�D�$�Q�;-��4nI���o�U�+K#A��%��A��D�alW#}W���[^+�5�;�KDa'�A~��5��׾��Z	�\;�6KP1#$"���>�[���'�������5M��v,�lG�;��`1N����F�a�:���E���;�b�>�.���#R���&-1��}AY"�������@Pg�p轿FF���)Tԋ}z����d�<�� /S��4p�v*��7�������)�կ|�9�'�X�ˆ�3���4��B:�5�F"�r��ܻv<��7������Ϭ.��ORt�r}���i�8���)��Ay䣃�v���:�ħ,$B�\�V�w�Kg^���j4a���p��D�!�`?u/6*n���!B��>A�!,��fؼD����)c�$�WJ��M��wr�^�$j���������w�X5JՎ������m>> V���|2�6���#f�i�kdO�w{�������˧d���za!_���~9�O�f���]l$�����F�S��e�/�i�cmy�hƾ_B|}C�l�������b�����m��/
�r�>����-�S��o����M�aA����Y1�k�x;6�ۮ?�J�]�`������n�=����S OEbORȁ��E�L�Ӝs�{��B��A@�
�Bx�B�:��1G���KXRɮ��\�g��Ad�R~v�qS�е�&E�-���Aܟ��ҞY�S�N�����(Ĥm.��?p�}gr�6D����H�ަp��- Q<|�ș�)�L�nenʺ�6<�c���d��j0��V}ņ���	Tᾪ����[��F�1�+�{��21�e��5^��OUO�D$�����-�����L���M�pc���M�W|t����K�_\�1�a	�:�#�Uq@v���28m��(�:�)2|��A��|V�G:`N���z/��l�7�]��+j��C=�
�2�l�i�j]��`S��Z��=��O��x-^�IdI���ҏ��ƕ陝	��dn�J������wr���b5uFp�t"5�Op���Lw�(����&���8�D����p���h�ͼ�����to�q���пs��cl�׮@��u��eaǰ�_�)� ��כ�Q�`B�#2p�����<�A\����+2,�8�u��P�g�0���=�_�]���a������d� ��HH�׆+{~⯡��˶���͒������;rBR~T`�"��*]h�*g ���	ft�|p�!k��+�w�Q��ݰ����,VAg{� �Ļە�%��ޕ�>:���NH�S�T5!���qs�_�D�[��n��A|�qla^�S%N�/q<~�� ����i�v����t�c�3�2a�&��jdzw��V�>�V[�'��2���x��j����9�"j���±9gW �l�i��>��q�a���.{�9S�Yw������ ����\^���ZX,�[�]��t�p�P�����e��35۠�M��4|L�	�L-83cQ�/�x�Y���n��A[���;�D]���š2���IH��4�n���h� �{Y@�9O�
�����FHsM�!��
�'�r(갵�JzF{rK��T���eeF���mVw��<�f��V�ժQ��0y�������!����Q8�X#