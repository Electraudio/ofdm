��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\Z^v���ݞ�ɜ�0�����l���ŭ[�΃��2CN���E�=�����WL�[Kn�r5w�)�#�g<��QyH��4��n٭��iٰ`~����݇++�*��<a�PGk���k_Fq��7�wE�XBp}Q�_�G�0n��	~���F��S�/Ȁ����ޕ��G�W"'j��Zڣ��dIyt�wY������P����b�n��R�+�Ła���[R�7_��i��`�>zSQ�ǥY��ف�ru�e������z�4ȸ�J�wW�%�3�;9}\o'a���r�,_ǁ�n�W�*����Y�sҪh$^	�CJUj���+Y{���/xOq����������`~�?��b)�`U��q)��ȸ��}�Yfj�	�Ҏ�v�q��'��ٞT�S��3ۇ�^�����fQ�Àaϧ�3F@R����r��L���ţ瑿�/d�4�T�]�٥A���bA�Q���x%���*6YiWp���Ԉ)t�Xd�FOɕAޝl�Ե�/�ą5&]/W8^ٴ$ ��D�����)q�A=�⼾	xr�f���,U�8e�M���l홦����lG�`t��	*�x�P~���a����5��;��`КW�j�J��E]�L	�t�1!;U������ȗl�~��P��>���n�a �<�9s�)4�w�"V�s�ȑ�w �lqŧ<����_�����K���$?��������:���-�_��H/�y_5�����в�&@���H~s��f-`�>��"5�L�v�O��u�Q`���l[�/'SE~�4����7�p��J;���Y�m}��:mzbGÒߩ-����4���l�p��	������˰�SJ~VU������,8�cV^l�.<8�p�s�_�:[ �K�YG�M��L�E0��a	nj�]g�׼}LE�~�I[�%4� К������ b����uU���O�y߰�l^��ϛA��	�D�"y_�����E��kZ���	��Hs��=�t�8�A���D����U�7�^WO�7Ѓ�빭5\��C�b���U����G�z�, 7�qb ����+�;��"���[�z7�K�X+t��O(�%��� �x�S�@��|($�����w6��OE��#����O^-V䰽i�	�(J����i͑q���$��90�����P_e��t�e����~�]�?�w�1�	:ɂ]
PG}���r��#�Ʉ\��'��mi���^[�{�aW�v>`2�K�O��NtC�$� E��v��0���x���T�%���J.�E��Փ�J���L��-Q.�<)p0�m#�uc.;ܦ(�s���p���Y�
Sv�ōA��ƍ��:Se1��i!�-� ��-��9�/�
���Q�8[8HH�N	p�d�k�̘�i����Nm?�^.Nݾ�?7-!��/��:e^��} ��.=����N����S��<ߦ_�2G�[m����R�\�t]m���*��]h�{�_�����{�夌G�?}	��Y2�������s�K\�뾛�pe�A�g"m^��"�t'�"̾�І;�K�?�{%#;eev����MT܎"���*�Ö�l,�R?��?�4�|�y��$�CQmC��D��;6F�j��5d6O+�.)I6��=������xփ�LeUpKk����F~C]�'����M2_�Xc �sH�d���Pw�!>P�Ƥ����j��6�3�+1:�g��'lr�z��n�,/5`���CsLgcU� �����i7��Gq�Eq�{�8vV��Lm��)0�
��a��"�H*�&A9�j���`$���U���8-�����*�4,Ӊ����+��L��;ұ�(B�o#����b���e���s!�]�i���s��(o%7w�V�O-c����D�4"�N�|����L�!s��������2cF�t9&�^���v���I�ND����f�e��*4��f��c���nvo�*)���v���S����C�!1]��Ǌ⚺�R'A�(-^�t0,�M��թ4ͬ�e@�4��p��Σ��jn+l��]U���@�Z��#��=fH�����47�)��G��'o�������P��	���o�#�n�WNl�μ��7^R=�q;}���Xg�0�lPTs�Aۄ<e��-1m���pV��I� �K�N!��+8��r���Zɷ�<�H���i��?�M�j��
)�����C��Qv��h���bՃ�r�:9Eq1?z�
Y�+ ��r����NS�4s���
�d�C��gP�׫�iioVVp����*���ÿ]�7�C�����Z�KH��2{_ %�H�8�WU��M
HpH�ʨ�8d!<��� ,왨��/0��-z�qo��m��~�4� �\&�C�ϑt ���0Z�Xڗ)W~!���+��^�t]��e�>����2��o~��Sҧ��w�L_0=��i�}�ʙ%/v�,�p@�_�zCf�so&��lv�vN���yޮv�#��)����3����Q���}����)g���/������s��g�������)I�L�D�ƙ�g�M��m-��	cF��_h]cLr��G������;6� ���s��e9���R�[J�����w�=nj*\�Uj��t;��~fM8P��%_�%e�6�5�6)����r�&��W�(�%8w،��v��H>3'�
��x����I��w���H$Xq�����aP�:�d>��2ռ�$�]�M3�d S9כd�
룶��b���v=8F���_]1��k������+�kY/��y�}��g��6�;���	�aY��5e�z�9gU��<ـ��/�1��e�ü�_Y(Rs�����KpC��X�j~ɷP���ͫC�Q)A���Mށ	��2��J��۫ ��W���H`�6�
5B*{o~�fg��p]0�����R�N
�3O�@S�`����8�3�ՆK���岔�W��b��C���XT��?bK÷<���>²�̉��TK��d��wc�Z�<E�W6^$��S���1��O{�֬��������:���#�$���ņ&kH��l�S^y��� .����!n��O�ĵs1���kt�*�G���f���'(j64b �+$z�ki16r�5'��{��O@��&�7hԆ�b޲��n���R1���|}�8���Y��V�fО��-����4S�c��G��WR<�f,��p��b9I ��$��!r_ـ�7�����e�3��9H���de\}��!�|��B<Y�݆�w��%W����$�L����4@���7���#
�H)����ß8ؽ�� H��<4`�[K�l���v��r�� ��j�=��j;Z�D�\��%_BQ<���"(���_Xkh����A�GP��Ʊw�a<D$����ˣ��>&��u�z�X� ��d�߽v���)I+��K��Y��t8�o$��-M'ԙ������.*�6Hr�u��Bt`"}�����1)�i7����Co��d�U������?\W�.>48A��`�.n#Ǫq3�#C�
�
�:��|_,�@)=u�|��{�I�t�\�a�o��,�̷Y�t�4�}���V�]t�pe���\m�w������M���}`>8�������S�"�Q�D�4�O�G{���t4.b:����A�v`��:�{I��n�c�8Z팖���/�fi�|<�t"����0��!�D����#�����C7���*Ȋ�M�9`�r��Q$����ȿ|w�!j#��?�"5�|	Υ���颩����Si��c�lO�$�~�4۽�E�b+%!nЪ�8��[H� ��G;1��k+l�N|�ʰ���iZ���^ՙ�K��X��SG��f�E��*�t�Xվ���&�U׎
94��3���`?�δ~!(@8}`J�c�(�gD?�,����/�k�9Q���CN��?�j��m���{I�����$3Y�����r�b�?F?k3|�7d��a�����F��B��9�̈́��AM��4����P�*�:WY@��0�928���'����4��oce�^�l#5g@K�;�/&�pv�6H�Lt��k�E��!� 18沋#���ѩ���F�wѺ��+ �B�/���Kq_E���o*u�a�����k����v��wӯA���"4�<v��X��Ƈ���	@A���e6��q~ń�G��~�((�e��?����ǁ��ޜ�I�^X#��Ɩ��~��� ���9Q&Mr!��*���Z���P�ΤrG�ܿ����AX &w�"�pc嗝U)����!͘����Dd�foK����m�Ϻ򟬚�t��|��尌d����,�4���|�r��|h<��AYE��jn���ؘG���$�ϟ��'��ҁY����Y~��J���Kcm�i����qJ%@�L��[E�k�F��޿.�X����F�4�ٷ���݂$G@9�ks��.:jѨ�xwB�+�
\W�`�9�1��3����ߜ��m��[��&��,���K拭������d��	�l��cZS���  E��-����~5�z��[b�	�s�,3�$lp\
Ig��+zct�$��m��uG�z2+aK�Y�t�Y韨��w�P~�jjmE�&�'4�V$ŏ�V�ϯ�޶E*�Lr�-�z�'Xcq�;ч��W
��h�k�'1e�,M��{L�;�� E���[j���$P(�H{50�k5*��\�Y�P�����jMm��F�w���tY�_�0G�8���G���y���\�l���M޲�d,m5�������ʹ�ڝZ O��w�wK8�2H�����؟�|AkCk̎3TN�'�\6�B�t��|�h�d[��/�7<p�D��ƠLi,�[t��_:�)�|��L�
���_j��n�ss��u{�"�Ru��P�3h����֖0G�������*f���]�aT�s���G԰��$�\_
�÷���i��N�
f=����2��B_N�~o�-��0�FzQ_V��Ț�zs��zF����؍�{N7��O@?Fʌx(��jD��AL+^����8������@�������o,�P�у���Yֲ8M�C�ӂ�J6W	W�e26�4��[�e=�؝*������_�C� �kb�i`�K�U���`�n�k�������˒�_g��uO�V��q_o��s��Dt���co��س;���
8_Z�Ѳ'/�@A�5�%���C̤X�'��im���`�)8g���[���������5ν��e�OX��j��#����I���;�%r?�)�i�;���((�>ه~@t'OOH�A�e`����ڛ�f��Ds�E݊<
	F�������O&}5E���6Y�ې���/��ϣ}>�)H�� _{��d��|��N&����ԓ�-��� Ʒ�R=v���b���(	q�K���mMǌ	�lF�ɲ̅|�t@�\E���]��Nճ��Kl�]�������YL/�´q��h���p�*L�-�?Z�r�!
�J^V
8S�$�`�q�c�˳�R�����6��I�y�S�;��T�(�_�a���U���U��8P]��+&l:!���~(�a��p��{A(�W}eT`T`b0�ob�����.	�H�imE��Y���UmpDDc�N�f6��l�ki�'9�_�ݱ���u�c' *_��e��P��&o%ӝ��m��uP��"�1ыm�{J�Џ Bgs�킎�skM���c��6����s�$Y"l�=�M;�н���nl�q�]�j��Q��g��DN�����U�~YG7��Re?�Y�a`zj��R�)�ϣ��N:T��Ef!>¦��|`��s�<��Ь4�2��Z��*���W7}N���P�^�)�۰'���;�֒�p[�	ML��zv�	_�G���g��PƄ�k��!4��k�q�94���N2�K;GS�1�}��/�zc�aS��Sa��2� ��6^��K�YS��{U�	2�
��;_F�
A	ۀ�S�g:oQ�E�)�TF�� ��glg{)���\��f;xu�� �=4f��%��PM%����
�O��E�]gV�twn���y�!�o�������¹�D��Z�a�'�G�T�^^��!�������L���録�����f1����|�k�n�{V+*�޷����N�兝Ȥ�G��$�_�Ďl@�q0E�V�Z$�0rgT���{�d��i����kσ�֡�PԐ��ފ(� 1S��~��Y$�J$����h�����z���(D0X|Ǣ��	�P���3m��agD�f������D�KL���I�t\�V����\k�{�� '&�
J�w��J���0fNS\O����yq�{<���J���gY�~���`N���l�u�P j�c#w�������r
/rR9�h�0p&j�]K�5H��H�� �O����)�0�W��5_�#�i�I��|C,����t��c���
q���#ɝ�X��CD����\>1�;�SS��.'��+E�\[���5'H��w��qnB�������uB��(��bN�$���[0�-t��!�-s�g�:� e�|��?�M��8��Wu�·��/��Z�n�d��͖�A�*�k���1��@��dZ���
�T;��}<�_tWŽ�	����.�@�gV���[��)ť�{�����@���ز�+����O�煎���^c3,K�A9(X��!�֎_�7�8x�y1���:��Zr%�bfk�Qx��{ղ�N��������"�esK�KF��H=ɘ�����fg��5�"�=�\y`ϲjJjKs��Bj��\(�i��W�2.���90KӁ�bw��h����ar^?S��$������'���!<��Ŭ觢�%A〱�nRS\����������*7t{��3����rE��VL�t�T�p���T;�7�S!p*���sI.�T���f@ŵC�R�S`��B�Uym�@w;�=�*^� ���Q+3_&��u�ݎ�Q8)����s�,)�
a
�;��x�X�m,<J]�����	��H�+%t��$@��L�����4�9oɢUm��A��q�U�E@��	���Ih)Y���;�Aຉ���Mp�"-��s�"=j�4<��~y�&$ȳ.�<~�L���}����fn�� *(�!J����W�Ђq��L)hngȑ�v�'-hu����O���Yi����b����R4�KY�[�Fö�$I�� �n	)hu
�9��|M*���8ۋ~= {14����}�|���d��꽃��߸�r�������r��JӮTȫ��j5}�.z�`�C�z<E&3�����s�W
�Mk6r3o?����Dd��zR�5�ǺA)��^��L��9�l�=؊�4�=]�3>p50 x�5@��kC���	�<��@$��RN/P��ww+l�A�s�Si�����ȶ�@Fe�Ruth�"r�� >4�M�=w��Rf��U��m�p�	+d�e[��'�\�Lʗv�E�O�VXa)��v�xnrl9=
�K�ڎά�ٓ� ����&;˟J��:��%�ȣ?HA����$#��-�#�}�У�@�&�U����m�([���9�ϏKvM9�c�F����˶ s��=��M3��ɩ2AY5�+4�|�ߨ2cj��q�"0Ȭ�G�T�i/���W��'���97xJ�ZA�N!���j᧵?
I���k����$�PAf��mګ�\_H �4��׿�v���Y�0�N�|r>u��wMږ��m<���$b��9��f��0DϾ�i�f��<X�6@��^�b��­���7=ʽ��:�KBr�sGWޓl�I":����R�D�t$�N�Y'�T~�I�X����6��H��.y�p�~	_N��~kJ�_}��g���ޚā߇���P��y<��3y����S2%$��IR��X�r� �-�����/�V8�y�k�y�p���C�
��r��/܌��}dM(�x���g�^�I@��z�>%����Wk�j���1u��4Ԡ:�hE���Ud����ݾ۵�+��p��ְ�A�0pvsL�(�V.?���	�z�u�L܂���d���+�k��[����Q�����G+RC��O���5F2�`��V�`t����av����u�ǔS�	tyd�+ޣU�v�žQ�����Qc���DG��&"���h���^m}ɣ�j���	 ��c�T�m&ı�O;v���uA R��
�Q4��7�	P�L��m��{ �Q�6���Y8q�k�x��ճ�]��6�d�IH��d�@8��_B��gӭ)����eu�GV���uR���JyỷұY�����!���B
���3��$��ę�iF����JgR� B��%��a�-�m��o2Lr�0���
C^���d"H���RJ{�)��k{�]��`X`D�t�d�?	���D�����d:S*zcO�� ��T�#�H�Q�R��4�)��f�G��1i���υ8�.�M���qm yn�>^a�W�f�{��E��+����u`n�y&ѹI�5,��U��-T������"�cS��������t�m ���D���F3�S�3�����Y�>�.���E��r���Y`�9�v��A�q]-��T�Z0"�J#���j���*�d��#]U���Ұ��ˊr1a�@����[�����Z�12�	�Z�D9�sƇ	G5�����N�<-����x�JkM���̄�4�svՊ��xm���.�Ǽ���q�y��Z��#�R���F��yd
��T�_[!Gz����2���M�A�#����/�uǈ������=��C��f�O��Dz�GM�<w��跅�g��l�����D x�Q��X��\a�~%��nΦ�(|=� �Y��,V�;�G��ئ�F�����at�����&��>X��4k=��|��c�)y�0�Mf����W)������w-��{_5ĴEw��{R�W�΋�ߊ?=��=l��ɤE4��`��z7*�3 I�5G�&Xv�ʱ�ܠUc��P�S0Y�+pߚ�|���l}�9.zM�.�M ��2'mq3��BFH����
H/ɓ��������%Z�3�t�RhZ��E�N@uIt��cš�J2^F��W���-�6м�,�����u)Yx	��-�	���2�	�4��Yld�����.�Z!��y]�ܚ�[?�\�\=a�����h�Qw���$Y'zrD�J�\ſѢ)�8A�@�BN0qј�-
�8n�N�ؚe�.r��ҧ��{t ���)��ګ_��6.ja�1�ϩ>5(*��aP�:�TH��$�jb������b֡��	�΁���',�RԠ!��%#��L��&y�O٨�KU5��m�k�q4SUT�:�ǣ�^$	���'5�#r����L�� �~��3G�"Ħ�B�v5 ��I|s�
�|R�\�IL�k�n��g`�=��D,����\��?�[�ە��ѻ�֨y {6�8B���(���5U���^�G���n���f�)jE�VGv�Ǜ0!y�A0O��N�{�Mu���0!�%MJU�dJO��Z~5����� �ú���x�\�����i�t�+5�k�|ã��o��`[��sܻ�q-���ߏ|Y'��<t:֞�4�Ǉ��Moj�-"܃������U��x	% �b�𲯗�(��i�i�b��I��!���'
~t� �1w;N�"���֞x��}Z��Y�L�mw}�ޥ��VI��BK��XYS��k�:�E�o����qV`~���G�V�{�)�xln��鐛jq����Z��yr9N=�oQ��k��io��d�5Pѹ(�����V��m�����?q��Y�V |��x���\�浣>%�v����U�ϴ�nL�������.d�Z�Z�	�y���1��K�J�x�G|��ng��Za<>��o�,�f#��L%��ߤ�\W�c{݉�ҙ9�h���SZ��XҼ� �l-�(Ws�6�Kl�dN����8C�S�Y�M�	��B�'����� V�W�lN=��nQ	�7��h4 s�n�Lc�ݤެ��\���e�ǭNv���;%w~\�ԥ����=����\��\���k ��s������{�����ONGt���q(���EeŁ�8d���8�tW�J�k��t�qX ��C��5�d����Z	�����k�T-0������L�W��Bōs�j�A���juL��İ��!<�)9���8W�65ȄpL�T�[�Y@���h�UN��>����C��}����%N.�%�2[~�4C�nnrhKC�T� ��4�Rۇ�V<���ð����6E��+�,'A�?6X*�`qO�}e��j���bā:v�KТXI��w2��͍͗p0FJ-x`�t��$�\�l�cb�`fF0�Fy���S|�V3c��Y�r�%��殥�a�����P7�� ��"��HH"j��t��NL5IC%�<��fΖN1Bw����z�H�ZV͹�����?̳W�|�3}��6��3��C�kE�H`��q�O���u�8�����4�3VsVӜ����l��?7	��-4��w�&{��b�ߺQ�Z���54n��8"	�Q�����b��=y,�r�;�/�����v��.n�$@�Oh���+��M�aZI��0b ~{�E�Y���:*��a���4l���0�*nW��Mb�+pM��59���Кr��^��Β[���c�w6���-P��v}�Ƿq��dS)�A�(��	����Y��`�B�9�Du�V�cG.����-��{-�(��c_�1��U�^H�St�!�"���,|@�,5���\��?b	�����2���:����-?}�D���q�4"j/ �{X�l������U8�"�ג�����Y�7��� ��������#�̷�W�34^#�W��Z�}��s�?.g���^J���p��3_*���͡�� E�+����m���N�eu_��	����֜���.��Ә� @Y<�r��)Y5T�2�m!*�=p�u������{yf�*Ȃ9'����P��z�:�'��m�k뮸}	Ci�qlⵇ�b���
��U���??\���u���]���7�ό�������B�-�R7b�@^ᛯuhc<f��
��;���5�P�ϫ������t'�,T9�qZq|n�jb�׶�l��IX���9.3t�ʯ����o+�mKM���d�H�S^%�R]h�5�l��7EZ��}���y�D��2�a�	6�z�+
�~8o��$���O^�q7gs�n�i9*�YaR[r��`����A���8�oNf�`;�\)��K�
y4}g.����&�Fg��ɉ���?v�Rj�V��ڽ����C���@�u��U��F�C��wx�K��SN2Us�����^:ϸ}+��eqŔ��	��k>ah\5TO$~̞Ղ��t^�ʖc��Xժ0d� <��W�mPt;�W��x�緃{
�}�$��8 9���s�i��n�H��d�y�_.C��9�<���!��.p0���:��,Dj�$�H#�\������I��tD
��g�\ ZS���k�A��#�e0F�"�Q�[����:]�{�%/����D�G��q����װ�,ǢA���qw��;�˱���R���L�R��HT��H�0�*?��G���{[� f��s���z-Jۤ�-N�^�e��(���i�|�zH�����;�IpR�o����T;d�:L�5�ݥ���OVեܗn��nvОw�PA��O`����]�% $8��؞��A�Gb����JS���˃��^�u�?���E��[!J�"���� |ԡ���a��Q ������ES��7�e�/+3P�y/��$����פp
<&ʻ��F#�%b�x�D�=54n[�ө��l�p:�ZMWZ�^�fG�gح���K�#�@�JK�*�ro�� �:t�r0���>�qG� �fĲ��ϸ��5cP�/�H�jZ.Y�9� j�D�SB_�T�`�_�BzZ�y�(�V�_4��N���q�͌�rW��|�T�`R����O�RS��(S5RT��%�Rs��|ǳ�V2����/3*�qT$���-�P��(�s��o������)w�����c�^yBg)��Z�Q����,�g1@eN1�0��K!��9��E2��$��>�%c��=rn@ވ%@�R��j]�{ZOb�����!n����'�S��Q�H�姘��k#��&*�q��S�^�&�0�[�xА%��j�@hPC�j��E@��h@G��ʗqǐ@��<�?��T�A�%���6�����ß���C6Lǉ��Q܆oZ:�4����|%�掜-PtN�'�x�l�_n�>^-�>e���F������f����=_Tph~j��R}���,L��2�s��]�]d�!AjJp:g�E���_�8����i���z�(|�1�/����Ľ�!����s*��T4��8��%��+i�ˈ�[V���K���)
���ǳ<k1]��5ә)�a/>H?#�'*kH}��f�ǂ����(���k�Ry�Hģ����u�!�Svg:��9X�K���V��R��?��O7�G�٫���oP�];�1�]�!�4���e��0�^����)~B����d�����	-Ę�+�������K��v���N���iuߨA%t>�%<ޞ��K�Rg�^���5�;_���N�����Za��6��;w�L��pW�
�,+���������0׶k0�h���P��n�;AX2mi���Y�?DG�r[{��%�6,������+Z�|V$=���(�"�*���ϻVϺ�U<<"����~t���<�;4Ou;+@�Đ�3�mT�hy&����R��ޡ@0�~}S�ˈ!�rg��z0�ҍ�t�ieK�`���0�ܧ���Y)g�(������j t��[�Y���:B�>��c��0�>=^@_���}&V�c�%�5�S�������6�bϓ�Qnȭ��3G!1�U*_��!T��ֶ�����Y��k�J�	QV�	�9)ir�T�O�ݽ�jZ�$�׃�qBo���bVXȐ�3� � ��䬷�%�(ܱ+�P�M ��YUgM}�E �~�(�S��%���S�(�%Ru[��K#�&j\�Άb�mC L �&���aB(e�;q���p��fF܇�vo�hr����ed&ۖ�ܳQ����wL�a?2�|�ٌ��ɀ�}u��H�yՂx���a��W�(�Er8��31t�=]��x�(�CQOM��d�Vu��؈��6	iP�d���~c��z�2 �?�Q���0����C!�ɦ5��M��f�?�vޅ��l���S� �c|I�~�Ѕ����������=���@:�g�\��]�;���#�!�(�gdP�E^��B�A��W��ߏ�%���==�ۛ��h����jOM���3xPB��#[̮E�_��j�[Vb�Z��	�ō;�nt����O,Ap�ܥ��	瑨n]�Kwٖ�4��W�1�H[Q--˘���ؗ���'8�tV4|���ʅ����}��S7@�
dg+�!LԆz���5 �/1��'��%����ʦ������!���"�	�A�T�?�O(�Crll�?\��2%�Vz�ݩ�{'K/LqD�������o7�w�h�^��7EW;B���C�KY ��AdMpVS�B�R׈{��|l��8�{N�W��C�2��EԹ�@�{�;���H�O��g�:6�`p�.�tL=��~r8`�m`�D��_F%�5z�����}[��u����Oլ
�[����t���㐥�Ey"-��+8�c��x碇��F	�2��`���sŗ��S��������W��6���QfzA �%��z4���9+�����o@@�PN2��Ȑb�M��%��x�L��J	b��!}|1YO�۝Z�U���~`{,��
�F9	��)E[��
��E�Y"��\�u���B~��  5q�?����l��@O۞��C��w����U����M�(�������޷W���}�e�s3��)�.@��ߺ�¯�.@=�6
�wh}�W���$�$G�MV����
�x��FbT�E�/@�-�����|H2�+�.A����ս9C�I��@�I}E�V���^T�_�ҋ ��V�\���A0�tJY��IО0��2��TJ9��*���D�c�,C�`_�ӡ�c����3���I��a�ܘvӬ��r��\8�C�Rj�O��S,��3��7?m͐�½K��	���Pʒ|�	����C ��f�r��._X�6��|�����Ţk��vSτN?��q��f �P��ԅ��/�3w�c����>:EO��=�3�<y�\�����W*}<��yU�����|�FP���Pt�g.$+��2Ka2i�0\'����a�I%+��y8MkM�H���?�_L���r��孭�h���T�~u��f��k��h=�v[} ��gW�B�a��W���c�<8g"�X�l-���`�""�O��i��,O��$J��2��3x-���r�)�[|��o+��E�$l����JGh�CU�$���E�Om����Ǵ��&#�-��<��v0��zQ�r����b-�ior�n�s��n���e�g^3r��1�#N���{�Vúќ��R̾P�[�����{�L���m嚭b���}�Z��T��w������(� �B���Ҍ8�]�8Kx�[E���݆ܤ$�	��r��6�@(}�C�W�ܤ��?lc�<m�y�旪���I���s4�v
!�(���9F�`|m6�rM��6���}\ŭR��J�m��k���R���s󺽪�nlN��z�S�@�� UF����C�=�D����,X��؅x\l&���	�������B��o��a��O���}]_6n�Rk[^|5n 2}�Șy6�'H���z3�fӎ�_D����	Ǻ�]k��v�S!K:+�Y���F-��J�#j�,)h#�a~��7����������K�c���zǿ+[oK���Kt�,,G5&�'��UF� ��n#Q�,K.���jq���6�8җ�50HIۋ�3� ����� 7���͌�@�e��;�Փ%�Q�
 $�(QA����S��64���V�����ϭ��N���䍥B�{�s�m��d�2�����SR���3��u�M��F�Wv���Pk��f.mV�Fz��F?���N�ܢ��)�����oʌ�M{N�B:;���5��ne݊.�����*Aa��0�b��͝��,�j�<T{�q�!ý$\O�䓠����m���!
��1����\������IK>סI��}����%.AbR�8\svp�	d�V�b�����0�Wg/9�ߪ���_ɥJ��9f}B0�����;o����+�R�,�F����4�^��r;5F.���Ӡ�<�	N��7����n@{�㟂5a�����#���ikE���<�����d.�	���.�����ochƇ35�����[,�n�+� 6x��d����}�?+?�V�FB��VUFP&�L	��⛴�$��!�c�Eo�k�U¯����$I�S7�t�ڇ�(�=ԟ�p�M�^\:N�٠�$�[q�z������1��^fu~��������H9�u<y���k�1��i�I�}��zCb�q���ڲea0��+��)q~�n4�@��ĭ�nE1�*�ࠣ�3MGO�-~Tf�B��5���������]�+��ɫ]�8��jKղ`R��/�f�g�1�ʧ(��6Ou|���T(;vr�Z7� �`�ί�"M���g=TLz��5�S�y8b�q]B�,D���5�#�#|dS%����`�q�b���KD*mMә�N��V�h\��6��c��BLo�0.���M)�SO�d�Y�|0e	��KpNLʼ�ߖ-����
�p�.F�A>�G�b��zn�Cn�m��҂P���ZfZ6~��zJ�mld
ܼ_��(�>��#���dĕ��('�r6o�]��=f0:t>���˄��	���5����������	�#m�9��������w�Ӈ�\�_���3�	C�u�ͩ�+�lg-�|f0��N��2l�U#@��T[ h����J�`���#�A�2�pD�O��iw�>,v/���&���3��:7Q����m�VTv]�{}�^(��[���\��a�$Y�ߗ.�G�ä+7
��B/�TI�If�_��j����wA�ސ�����CaJo���Z��amU��L/re��@��ȷ��K�"��:�,X
��]^kGA�0 z1�4�Os�֥����-Y���l��� %}����V8�{�ڔ��(o�'�x����WX�R�Ƨ�H�st��̋k��U�/�Tw���&�s@<P���e�0�.O��6�.�+�i����^��ǔ�����D��&nU��_�y�.v�mۚ������B�[��)�������l>!W���kڸ�ꤪ�e�� �Y_m��҆�jC5т�4��:���#&���:>o�Mp�עϨ��j�$�+Ҳ�0�G�\�I�sQv�	��X� 1S_cG�9]���U�i�տ�������`'�읂����L�6HB��^�W���e/|��� �*��A�B���$�S�\���.��O��/��Y�Zn��u-<�=��͍���ݪu�M9w���Ý�N-0/C߯$�e �hnH*�w]��R�`o�?��Q��H��#��>k(W<��6��GR�=����h0�E��<��n�w�2�k�ʧ�2��t5����,"f�Хg�	:���ܣ�5���w7�G
�wdC� ]�����Gxtw��ݐ�Gv�&�8��B\�5�Bvxgڢ�t=�1�;���ޅ�c���X�P�6zڽ;�k���;��[mN'�� Ձ}��S�nW�/��Y�3_lnd�+K�#�'����r�X 6Xß0���9����������n��\{o��r��4'�-���a�5o/c�H<���Yv]��������/��
3.�t�^�N�w�tv����j��|s�p',�);f
&��k�:9p��Ϭ�^�Ծ4>�R�/��k�D�B�*pӏ�π�Y� R�J����K7 HbO����Z�'O!�(
��x�z�]��y�Ǝ�!X��e��}������Df�
���"����n}�-��s�<���~tP�4:�B�P�F�Yz|�E 8�ņɅRZ&���ˍ���EJë;��B�\t)�/¦�/0���X9.s9(P�1o+ҜI�K����QŨ3��)g꽫����=p�P�͢��&�IE���H��7�+�cb(�Pk�2vb������E'�ҋ���k^@��!�G��`�
V�duN'Z�MĞBe^���-dX�k$k�oI��8��6�t3�d�(<0��C8"3�r�0�O�[����`뚺P�Zy�Kv�aZ�	�x�7�4�-�\5�*ߵn��y
��8kY��#Jw̴
�gX#C]���5/ۯ���Ԧb�:p��RMf��sk\�ї��;��l��� ׃錵�.�ɪ+�/�~j�b^m���)���>�zc	��Z䠜>=8��Uq�rK��cZ�1��h�S��ȕi�bi:�qt["���%���u��3�ZЗY�4�ͼ�sR؝7�B����%������B��6�er�d8.u_�Y��"����t̕�"�]z��$GLq����9�
]&?x������wLA�^�7T(�" �?@��1�ړ��u� �`9�,��r��0Ҵ^���[�m��jؙe,�wV��	�v|�پ W��ς�Ҕ�p���t�k��7�=-o�L0�F�nF_!d�F�"u�A0v�"��Zר��Uc�[̠�|���U���~��0�P��M'� _�k�L����&3[���q뀖���tR�A��4Tl��gP���VOO��!��!a�~��o��:_���I��g�K1��G�'�5���)�s^�'�9T-���&S�ȉ��/`�I���eL����BE7]�|2��"�������l����OH8	�H��E�]=�QT��
"���Ʃ�O�۽�G)4��MZ)y�SwzXхo���M��u�j3�1V�\���#�w��X��9�=�j�v4�����:M:��G0���h��� 64�WC��3���z����	V���9�P�z�v��"s�,
�� ���bX��S�kTH�+��a���8^\t��7���{����	�ǰ��VR����7*�ݠ���X��=bf$ƛ�'����s�o�P4���%�7�����hr�����N�nv��!a�!<x���B��<�<�!����v:�$�Z�+��T�O�� X���[vX>n̼'|����n±��b�څ�nɃn�FQ[��p�7���u9��$m�:!@�5��L�s�}�A�*��E%����S�tH�Oڜ�(����f�!sC���4V�NG����J>K#�Ҧ��Q=�SJ5=���FnS���N�@��yH�Iv�=}�PV�C�:��qu_j"�jl	L(03��.��$�fh�?�k��m����,"�����*���<�SQx�e�,KFF�rkr���{I����1�^�k�5c
E���Y8I�K��A������Ω`��~���F{B6a*�Ϭ�~����j2��*�>>� ��s��.��:�	��uj�������u0/�)�<#�.6a?����*��CA��1�ʾmUx�����8��.	o�՛zԛ���	�	�j^�]zu�'W=�8��Z�?��B���;�0���Ec��X>�\R������r��;����9�Z5؅8z'�5���\��8��ŗtz�Ќ��1f�g�{_n�U��5�?H)e3�+�Y匥�ՙ�F����2=1ʘ%vu[�x�Y��`���dQ1!t��c��7'I(8��G�3h�g�Û�X5��<p����́ʋ�;��~u^�<���Qh|>^��Z��a\q�9�5Z���YY6���Z<>X�p�H@0f~F[W �c̢��J�0�-�!��DZ���N5���{��u�8����	�]�S����msaȽP�B�l�ױ8�o-�n��g庣a��{�k#�E�%����G�~@��3�w�&7�:�	zg	U��&�n���'��떚~��Ř>���R8�S�f�&�r��Z� �_�7gB�g�K�U�Ђ��h���.A��z������[U*�v�-�'`U��:ȍXjm��ؠ�c���
<�=�r�+�������~1%g���O��qrO�@�v����{��@n0���[�:9����hK�n&�W��|h�7,�Y�ע�vg��?���L�YUZ���`�	�b`Z�r!� �G�˗JO!L'2c�C�����ޠT8�#�͊R�b�~��l�^RT�AM���U���3�R�������e�ڠ�ʟW��Cq�9Į�o՗�/�ӢK�S���ܱ���5�+�azs�&Q��V�^X+`�!
�x�x\�d�ɛ�(U�;���l�EF�C�pb���/�w�YR�͗X�T�"g�	�y�NR����߰�˪���W�E);sN��Q��%fE%D>�H������Q�y#��"���ŧ7��j�ϯG(6�z���z9?J(�Q��a.�G��#��V��j@)213ZW#jY�| )ɮ��}�!*pDՍq#A�wy�4�s:�����;��u�8�&u�c
K�~ޙ���A.9����}��B�UΦ/�@�cV�B���'\�y���!� ���A�b7b5"d��С��^%��#)�W��^����d�3?�e-~Zu�W� 
@�f�]���-(
d�E����䭫ӑ훬He�UZ�'#I����Ë[�j׷m�������"���4cUܯ���g4�D�����z�^��jY[u���+�k�>ϫ���:� 깉)�7��RGK�=�@��ʇ�l d@��g���� 0����Hɂ5n��+�_��~3� �2�l���g�J��.R}G�l�� ��5/���C w�&]E;�bK���rҝ�k>&Y��"u��#����4�7�=ܖ�?^I���q��"�Ɲ�����$_��B���j�������������K��Ƌ\����.��W�T��Ɗ>D~����q��չ�6�-�mRưl��& �=������/�L�}�5��l�4qh�!:�L��z�'U��������C�Rc�~�=<uFK,�KّJ��C=��׳}Nk]��U��c��^�a��d�j�J\w:�ɄV{�ЯZ����� �J�v�-��-�1{Ў�4�1��}��HL�0��B$c��^�*������U���`�4>{L�3`ҿ��Z�B�۞��KSXɄu�L��CT��t~�-�=>�g����(TdO��<����[�5�T kų�V�+hZ�,d�(�l�"��v�.A&8�j\�.sD)��ǽR�-�TM�
dp�^X�`��3�k��0D��5�3 o���Qi�(߅>X�+�Mt�KE �5��Z�����G#.``���м��%o���.�_&G�[�<��?��pS����=��Xo7�R޽��fO�Ka��c}�2��[�jD��c:m&�}"�jЙ�Z��0b=�a/����p�����Qp�>w|'�"v���>��[�x�jV7w����F��XC���r��&�ٝ.G��� o$�vo���Jt�G`��h��`��3j/C�tJO8-P�%%�p�׍���z8GE����rKb��1ri��9HȪ������!�N����3X#!p�������9��_My�u$eH>�Z|R�6��be8,j�@0�b�'�O}8�锝i�T$��G(�π�J�qx�Ռ��G�D�>Z	HDSK����n�svW��?N���p��*��y���h���s8�����@w8���<{z"�E�.�<>�c�Ba�|�|�ݛ~��5@��W����@�jˎ�6�@`����4���i9���:)�U&� n6�N��#ʙ�>7�ec�1����޹i�M1GE�K����@���b鮥�v:$
̞�(���wU��+�Q�9K�¤2rA���W��u�!�f
�9b�ȋ���Y�������(A���.�:R���:UH":��u�Y�,}p�v�8��8kqH��u+jA�Y6��nG�s���*Ί��8�Э �~aܖ}�֐��Ĥr%�Wd��F�<��̼�K%W���ΕB��(�7 ?��I���K�',0,ķ<�x5ǟ��nMߛV�O�P\
�^��/D��z�/�%������*�Қeh��D	� ���x�S���V��k5���M��{��и�y�Sk�[�&N/�ӱ��vOO��OP�V�>��J���g��RWɣQu�n���j�d�A�-��*�M �D6PD�"�e1�U�gR��l#�]=9w?��R&߂����@���&h��TG.���V�IӃ�?\Y��e���Y �7l/��Q�wsK�6mc�̲�s7�i����!Y[4i,�ϑ����#�g0��v�;��I%�Z��Y�x��j^�������[B���N]>�	D�#љLfԀ�S7[����A�G������$�A4���#�/��˞>X�`�r����P��B��#u���JBV��0�QK��/��a׹�����'�W)S;�C���?�y��.~"˽(!����q6Z�;�` �B,yěE��bAT�*W�;��@���0#�;�{ױ��s�2��xY]T-3��x��F����f�k��2����Lr�S�S��6��8+/BcP˙f��X2�zV{U�f���K�]�Ot0��t�@�͑���Ur�O�Z��bǶt�*�/��K�}�[D�ꙩ�5ܷ����H���fS�c�@vgD�9C2e�ք��~�!Aw�ړ:����W�a�$��]�e��y���+ƌ�u}Ntn�b��o�S�l��/SVw�_�ݶ�譖E�: �	:p�,Mm�6-�t1H|�A�3�%u}Ux�|�?����~���!�-��ʦ9� 1���з�z��-\�o��載����BB�65���-̝#�6�,�u����U �5Ü�?�Ql�eiZ����*�/�%�ؓ]B� d$���:D��ZV�]���lt�F;q��d�C���=� ��p<��]���L��q�,����!�����	5