��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^7/\�ǘ������W��O[b�^��nJ������`Zu�i�[��Eu%F>�,��ry��� �]�U� D!� `{�RK�ф�9&��nZF���(s�w��x��ѯ#�V�D�D������]ӵg�d��j�\ �X���SBN�?�&��~�o=i���	��n�����«��>Y�7�]Y���ǾW�S�H�������'qs�+{m��-��7PE�=���D��3Y��po!呻�-�T�\"�����K6���OMŦ��G�$��_C�p��%) I6� +k���k$�ϫ�ס�κI�~'5*�/�'���Qǘ���6������|@��[R����.;e$N�VݩtV{-֎�E۸�7����T�2[�-�7qN~S/Ѵ{����=��=���ђ��;k����$ڦa��D�Z�,�����4D�+Wv�4-,>PhR��������P=���$�#O�� ����&��mTm5/���稰>di��[b�������.c@_p��x�`	���d�;�uP��e�J�1dgĐ0�_��+K������.b���w�o[��<�v5_�*�!�mA%�2�F�~	B���a�a.y�*�c���ܡ�m0Zs���8��k�h]6s^�Kk��;�� ���y�!{?�ﳡ���xk�8���k4<��owdo�w�����%�!��afc��f�H�oP�X���p@j�,y������T���*0�"��8�8��2E�ۆt^����oj����y<���/
�ym?V`E���eq�L��m�b���/��q=z��jO{���t�sG)�A�a�)3Aeu�u�pq~s�8�=�T,ך� ِ��Y��(4�?9�pouv����{�Kv�?�<��72禲����y�� ��ZI?[r5���"o���1d�h�<�R_��	s-���Я�����N�E\[z�hwW�*���3�qx��J@��*	��% ��7Ը�����KA�a��Ր�u���G�π6~Ng������_i��%���S�]dHw0�$|�XP�j�&$�"Qe����� +}5�!M
������?Ħ��t�q�Yx=�9վ}477Jި����"�����х����^���.mQ�?��R}��?#�����xv�Yťl��V�g��]_*��\�Wj7��m̔?�����{��k~��j0��޵ ���#N���ǒXLI�l��_��d�z����yٺ:��U��i���L;pvSo\R2!nE�=��,�SJS�JtR�>YɾE��*�����6+/8�+\))޸���:�������7T-��-�t�R(�p,G��
E����2�{�����ocJ9���=w��|��*�$)�As��4�f��+e�U�hG�\��thN�qb"8�ktrdժ���YnNx᪱�1\�r������%��c1±�h��X�R[�]�m��wy�!����������_�Mз��.����߂,.���;���e�)�>%:gϟ��Q���nz�GH~�(� .�˘�Q�ʙ�mg� aάH+\�cV�L˚_%��(�?e��=5����vgc���+��h-�cN���	8f��r��U��"����n���fZ�>�C����'��J���TxZF'I�4��YlkP���2�g��C�,6 g�6�|���O��X�ޗY4	�A�':��/���X'/�������VL!g������'���n�5ɛ>�w��g�b��'ף���TA��e6�P.O��%�U�ho����6�}kצ�Qo�w��;W��Lk�R�(�䛾k�u�l�����1\"	;��/m�e���Y�1���>D�����֒>p���X�	���vٓ� H�MdV�+���m��B�׸�;i�Dd<!��h
�l�aM�&�jD��F4�/�~�h����R�\(���[�H�#4�R�&t�5赧�ˮPf�H�.�G��ޘ(@�_ �����<~G	�H�Fe�V4��ܩjLnGP�$W�	�U^ܧ�2d��� v����q�u����6&^��fbU�󒌑0Q�����=�#[6M.H�I�o�O�0W0Ǣ	A�n��7����Iil��wsnے�l�f�쀐�oIȓ5t�z�ӥ�X��2v����}��[��ߓ2g��w*�Z�
*���:M��3c{�I6�]�9�I�R$
�%l�o��5�`�Bޓ]��T�b�������W4�P6+�������Ȕ��3�t��U��1+cc�]sDךi�X�욂��ud��O��PGyu)�ߺ+W���\�&��_'@���!~��K�"s���y��*�&����r���c�1jX5�\b�b��/-P��Q�V�ka:A�$�F [���^��s:�3$;f�/�jW�%n� ��;{�8�c�2:�}��BU� �a��ת0�e�2�A�K@�SN4����c�Q��~���5��o6܉�@�W[���_�m�2Q�����6�e�jZ�cZ~�h�V��ì��O��^:�e	�A	�����>�z�1�J�W/��t�6�j;C�5�@B��#�
l�XD]�Ǖu.����ޠN��iIm!������"[��-����u\�׻:�*Ԝ<�/rW���V�O�V��Mt��VM)�դ�yq�C���e֝����6��8.����6�� 
A�;!��iE�*��+��m���P�\��K�!dc�1�Ӷ�q��fЍs#A�7VjL��p�'�i ���������,9qQ*K[��_���PT�&��(K����B&�Ȱ�;d�7}���y�*��U2�9a>���ƥ�$�B�\�2��#{�g�w  �e2�n!e��$7��o��� ����
U+ڠG�9i���6��a12�l�7���`,Y��j����&������ѭ�*9�e�/��F%Z�ޜ�5���d�8�P�VxF�>�`�'��"�E�4l�à�HsD�z�t���RK*e�	C� 5vA�A�1�j�H�}��}0LĿJ4����j�
U���8��b� tѡ��q��S�k^%o��5�\QK��$`D�*�y�o�u�[��t�Wʕ�L+�PL�M�sZ�{��\3@v��o��$�&��0�����0T��e2�z��7�H>��9�Q�����U9��/J�ڈ-�jE�O�ǅ��rT�
$L���1�o��*1���DÍ��
��!{
��n|7}ћ��PhI��#�#����r��X�����A��c�I��k�@)���_�Xj�t�16>`j3i����_VX���h�6����h%�s�;�7�
�K��������?M#��[>�/(b���M�4����9_x%tR�	�k>C(e�Ί�1p!��C"A~x:MP�k�m���,������of\'����X����  Ц<6Vi�W���b �����dۧso�#�/��D�4���|�X���#�+��H,E&хO}k8��T���}���Q�o�FA����8��/[�-7N|�;��1V�C�q-y��<�K	����DP��:LƫY���n�D伇�ś7QF�����k�Q&��b��J}�<]�qg��O?V��^��}^.F>'�wq�&た���o�������C����蔁y'X�w5���=��>��'�Y�����/�E J3֦�3��fPzw��5l�׍3=����آ�����K�@�e��A	��8�@��;��M�y��1Ģ�:�ũ���Hhn�Y U�/�x<5� ��U�-K�P�-�n*|��<)�μN�JՔ���؏�/�Q;p[>k|����ݦ�����R�z�ߗ;q4),�`�$±n�H�_�V��E���Z�����]<���r�G^���.�6��aj���M��H8S�CU?���㙾Y���)��1t
N�?qUsJ�5����|Kf���!�97�aTR����`�����4z��whn��h��Q���nҘ�:\�>WC�m��T�LI�<|/  *C�O�<�!�ƍ�-��Ł�;	v�w�[��}2b"��z��8��&z��������9v��б�A��7p?�o�Pid�>��[����8��jy@�gQFw�+�40.鵻Ű����x8����\~�Ԟ��ф��r��.��'p��~ �Aqb�j�Wa�*G8��$����5*ﶨ�e\ۓsy����'H�TR��q�Uw�:q$P�te��/���S�C��2|x�h��1��t~y���@�B{$@,�t0@h*^�]����8j���\��Dq���׃���W|�t���.﹟M
�U���82�W�$N��ߕ��Ag-bz��P��yJ}0h$J����+
E�=;���L���A4�\"e�<�m���;���]Ş�>��|{(�p�zV�]G��|ܬ�EnDXߛg���i=��&�Ӊ��,��b�$����W�Л&߱�o�@Z��|z�C�Z��(������fyD�^r}��yV�N0D�g�K	�cݶ�l7&��&:`3	�y����2���n� �>�7Bp��� SǮ���dS_@#��,MO ֜'t ���a‫V8q# �.�;~s ,�u�O�1�?lK̩��[F�/��y��L��3̍�.�n]j ��A:vP�z�8¨A�.�q�ˆr��x|_�����Y��d�,i� 1R���m�x-�ÇO�pok�!P4�xPG��LW�j5��MEC8�
�u�^�t���E@/$)�(��8����i���&5�@!�o,@ߛ�%�����vy|��h�'�hi�	
�/��^�V��R���.;✯��jyV*pk���FJu.ى�I�>��� �s�(/M� rts�k�5'6o"�4Ď�GT弙p�{ke�`��6�\�mę�9���n ���#$�7����#�!�Tt�Q��L�F�Hu��2!��!�7�>|������~�:��pbû<��i���_��(nNC�hm誓]n�E���H]vV�-��\��<�s�D�)���1W�W����R�|IOaP8^���|湿�v��:��x�BDƌ:A&�	� �k��;����}M�"�Pɞ���e8���?	i��|Ԟ��t�p),D�YzJ��.��r���6���C����H1`�d+�#V�nܖg�a�6f��+��f�����2�`�$��MZ%7�Lw� �s�wk�;�J�!x�a�2�����l�B�QԨ"���H"��l�<�,�\D<^�M�UE�|����E@�N�{�V�;}�������)�V���r<�Z��>a�?I����LR;��)�ʇ*0��r'Z	�:/0�O�1�p�7U'���k��Er�'q~��9�tɂć�#�2u�<���%�M ��p9Ӯ`�'��ڢ&��h�.Ql�Yή:�<Cĺ�(?M'��ȣ��u�K�0J�d=���!g����@����O�w�R	��:ltB�5kgN,Z����)Ԡ�7=�M�w����;xZ�U�B'�����R��Q/Sv�u)�~�Ç��сl�&v�D��*��X�;h��bH' ���$C����������C (���A�7��J��l��I���u�����,���ZUgs��oUf���Y�ZF:4Ԫ&��"�����O1l9���{|9l�A��4G#ìJ�^�i���UQ�~�4��x-t���w	b1�r��N���K�?�Ю`�9��=��4��<�$�2PG�d��
=�p���o���{H��/�S�p�Z~GN�����1AFW�����]������SԸ���\W���$��v
�L%<s��`����D��+Ȟ��f�M�'V�s��~J�f���ޞ�=%��%4����R����sX���L5�a7Jq���h�q<N�=����
$�T���K��Z*V-<m�\$��H"���g j�)�^7%�Ť�	�u{���3��n�*����j�6�
Ǐ.��^��F4����`σ�E�h�y���I!�Mc��X0�%5	�����7A�Y�
�.�dV�k�L�]�a�,�E�b�DӟC����"K�x�cD�#�6��E/0�+%;���)+�/�ljޚ���6D'Q%/hd@�k��=�x�Mrs6a	-{q\�OQCi5��0�{�O����4L�V�"쫜D�H"���ߥbIP1��;n�e�I�q�[��QZ��C��w_���q�4��,��x���Ծ	x�S�쭶,�����6v�F޵	��)f![���lr?*����{b\�$>���	�$�GY�FCs��ك^^3yBp��{�#Ks#��I��5(Q��Q�50kM�ق;�{<N��y�%k�¤���0�R�����V�_��ҳ_'�g������l9Lc�N�M~$�F�Hc�7��oi"��Z��{<g�7��d�q��XŌ"��k�$��̴B�+��o�*��$w�9U�40x�2�뾹����7�PC���I* � ��B���2d93�j�9�8�����lG�V=S3�uϞ�~��H�U}fhw��L�L;n)
�)'�>^Cۀ�� �5�:�o�!Ss%�m�A�eh�����߳T]@B�<��k�?K��J��~E���@����HִA72(F�z�z2T�R�s6����(XW#��k���{܃h�dj�
���Ka�*��\Bsj�e��Xk� x]�~�?i��JP���9 K)�~\G�z��`� }�ݣk{i��ɄKs�݇ir��~җ.��z�ó6�Az>Q�b�ߞ��D�J9
J����=�!LM��T���Җ��GYPP �������Tao�e�������j��X ��A�%-ְ
B8N�)6}E����+q CR�:�̿��~�ztD��6teդm�c��l��v�,f(F?��nv]kJ�Ɂ��ڕ3���t��a.-�����xnc�p �;�l0���<�Q6�x�Gx�Ȃ.��o]�x���|�����K(=|a�<� ���eϫ�z�fһ[+�W��*e��/cU+�*�J��K�-	oN.8-9�tѦ�@Y�����\h['7�4A���˪���g~|��S��O��F
��c�z'z@�Ŏ�&����+�������%��$�`�	y!%1@���:1�)43q�K�cE��I�z�����@�s�M�����9E���$��Y�^]C��W-I��|�&g1�����]��׊�����g���pn�B�Giz�y������>g�o�p?3_�h+5G������$�#�����2�<�GD�����3q��ZmJ�w��:K��s�Qji#<�q 0[��6WFNt�����aʷ�V3�q$N�+����1�G�a��5X��Rv�=��T��9�c�fǬ$Zg��R���X��0���=N���(*�
���Z�fL�2,��ˇF�^�����P�O9����	+e��[��J2:�I�q�f� �Q��n�'�
ҡGf�l�h����4���>j�y��UW���H�Ɍi�p.)�[���A�W�Gq�} ,=��x���o��=f-��^;	G�U�9���W0tu�ކil���tX�:��Z��K ��P�da�i���d@(���x�¥=؇��$ nXsdue��Jņ���C<$<=�p����������Y����0/Q*z�6��5t��8�6�\�`��Q�~2�ה��%m-n�� �Q^�KQu����4A�%�z���{�+s:��W�F�f* Š��K�W/�ڭ^A����&|�z}�I�z
������؀sW�[���-7��pMG�#����S��d�Ǖ��:Ǵ�Z�%/$�gp��+i+=�����~�J�� �m)�Μ5�,,�I��.��:���нy��h�����|fE,��XUg]f9�-k����ߒ����V�W�ν��{䧉l�@�8s/i҄�q���(�,%���O��r�rBF�b�r���$B+W�l�:��t���J),��ذ�Iߒ��(w@m&9O��;Y��>	t���жo -ӜK�e��QqZ�;��ƶ�"��&�������O=΄��36�ٲ>�mY$ܽSH����y�	5�V#����[Y�O�
���> �OD��:˳��#�G䘤���I~�����T`�T�񱦚?c����"��n�]hW��I�-������^)6,�| P*7�����UE�+�o�n���RGo7s�1��7��e�Pt}?r�8��8�q�J�NF�@��,U��.��8C�!�a"����y�uf}�U)R�$��GE,��F�Zw�,݆j��o�qE�����o����P��-��m�H����!��2���첚1Q`:�@����wl�"Z7*���eg���e8-�9��~��*�Z���J+	}����x��&�Q ��g����(G�&!J�d�=s��,�)*TX�d��Y��m+e�I5�K��·�3��E&�2�l�6�����Hިx��6��������+7Oo�=���{f�X��{񳖂y�^`Ke:��a	eL3꬟���ƍ&_���ѸC�͐�r��p��9P��F\�V�$��㩓)��S�gib j�,i��*�Us2_��[��1[�����O�B/�� ��"�b݆�adO��+�d�t6[����LЍ��v� ��Umy�w�g��Lm�x��a/ ��tz�x�:^�v<��#ʳO��ы5�ElK�ѵ��g��&X�ʦ��:��l�y�G!��m�l�|Q��*1
�y ��?<ϓ{7d�m�J�u�w�ȩS�� 6�_Z��Nx�Q�E�����sZ<� ˤ۩o�υ��ب�A	�'t����K��(4I􄹎n�{�w��/��[��T����-q����	$*�\�[Ff��_�W��}օA1�3�z�#�\�fx�e������q��*��;ğd>�����Ǿ��;v�8�2!\nL_u�C�m��3}(�8�����WvJL� ����ͻ�����A�*{:��
�����	fE�J�ߡoSy��՘���ڢ��$�Q]s��Y]��C�F!M��A~~�㼥�o몠����i%&�RVӁ�O*�J��4�����7��7�*�كd*��} �(���V��A�͡)j�|��p�Y��0/t�˩�"_�k��.S��fҼ�
]��]�]��F�O|  j�j����`�_���"jW���i�D����/;���2�c���@����]���ɵ��إ�+L��)c�=�D��~U+�������e~Q��]������h�U$��R(���˭u'Y�&/�"�s���_��9Ŷ����}󫢯�Z�[χ�,�"�u)���N¡-)�����p��}�	�~!r ���9�Q���(��T��=k:�<���h�_ͺ{�W��ã�N�wG5-ק�O�1��/.e��E~A�S��ȝ�/Q_:��#�:��}�Yv�P���+���ԉ�̱�2*�x���1Wt"y��$gM4��ŝ�d[������8�#���b�aA$�O[o���`�����$���?W9L���ذ��^�$�'�d���<�<���I@fD�}�\:&��[����#Ԋ!�d�+:T�|�E�\�+|.Yw���^@�d�G�|��t,����2p���
�ڤ���F],��-��&���@���ϛU�&!ѰtK�vm<w��$��f	��L���a��Q��c਒f�\��Y��=� ̀z�:[�׋g���tI�,H�,P4�S��O�A�t�h�CI庨cQ0݉��ݧ���(���t_{��i�!
�o�-� �4���鋼��4������BL"��f|KԡH����b���q'dϭ_��������,#^:<�p�	�����>���e�+�B����)�H���I��@�/:IK^��(�"QADW�`$�����q̦�]}�AB��+gD>�I��hZ�=EF�3j���i�&����l���P��Y��x��;dv���Q��=�Lj�:ҟ�]���m٧{^YM?ǐ�*�)�H��y5�W#�nr<KSب@����]}9�REJ=�"���e��hXD��~�*�RK!�i�TA?���m���I�J�j��0�Ar��_S%���0c�̒��/ ;IT��s�����d����#��+�!0��:c�ƣ�"�Z��ir{F���'S���_Đ}��K��S�F��sVt�91�_;����8֬Ul�=n��5��-z����\��.�k����n�����3�҃{2'�K�� '�?����"��䄶�4ٿr����Ȱ���@��H��f"�9i����3O/�uD�Qg�"�(�O��-�î@3���v#�n��P���}���7�Bm�t+� v$��<�i�qk�s�m�h�S(8O�º��zUd�v+V��P�{��w�+*(��D�_�хND�ʀ�.ٓ�U8�����G���zC��wsF���h�)��~�FP�f����?Sx���H��9<I^O�Ek�-��^����W�`��H��cZWDޮ�{��$����G�(�!�6�Zb�tێ�}�V��jO���V Yc�#����~���ßFg\x�����K�ר�rH�۶<x GH�`\i�#�#j�_:C�~�HYg�h��P6��M����;~<X�=�c�DIb�C�+w=���dO%H�t� V�ٷ͋��!��&Z����g���z��Ĳ/��@�'�^(s����?��]���Q�G���F�	��L���&=�Ԓq@�+���wj�V���Pɴ$�{�7i�E�$��x_F���J��l�rZ�T8quΑ���x��Z�&_��9�OAyM�j��3(�J"�� �tOB�W�24k�yY �u ���8Y[ \9�N�ז�|vI����Isvr��b�9Þ��A�h�*S�� �s�m�UOQx9+XPbZ�XK����g���M��.m� l�$[�cB�P�����B7����k^C�/�G���a���
��� ��e_���F�����{�,Q��=�~���q�5�z�>ǘ�5�����T�Tܠ�Yu�s�*�2�*T��g*�cȅW_F#�p�}Է{���`�2�A��	Ȃ�u�J���Q����k�O�>ݝ�1Ȩ�ĩIj3-[27�ǮGl��-���,iw�0��E�L6[�J�gW:`��Z����ę���3R��~��l1EG�>J�J@�P���+|�xծ�u)�p<��)�uTA�?a�Z{��{��"�/���\��~و���k�.���{�T6ȟ�N�I��k��B�x�S�u��9��Yz��U�5�]܄�'���-��2?�E��)�!.FT-8^�B�I��H�c��JB�����cc��.�n�4�������t2W�ȅ$��X�M���Qc�-|9gޕZ�4�>	ćn��ћ�M�-�����/G�ς'�Z��85R��!~��⣍0W���xpR���&�$R��tY̽�<F�J�/�����r��I�=��E��t}�`skv!:
ʫ�-5Bs�t#�ס0���dr��lI�Ǆ��ʺҝu
B��m����R�����Ύ��pZ��`��Ã��2y����ߪ�$��|A��W6}ߨ�TΓ�&��t�C�Eo��o�D�@��oc��Й~�{;p�g8s�����x&ZY����a��v���x}���,+J&�!Cg�:������ʧ�������/��fH��ev�3	��X-�F䈠©��ŞfS��^��^�d �,�ڭ�! Ȳ9���(\�R�7dtF�Ⱥ	��bN�L��}�w�Ɍ����'����/e�٠��.�|79݀�x��dP,†� �CC�m�B[`x��^/S�9�SdW�8�����?�m:�4�)<�8�H�a=̚߸!��!%�U��B?J �I�ˠ4�	�'�c��so�l�Ԟ�<�9Y�$#m+b�X�W��W�]�K*�B��ɠ�9��O��&��C6�ofM�cd����Z�X��U�	�n��n;p�z���ә�J@#���K�� �]���GQ?�]5(5��,f�q
*��c��8�u��EE���3#�]�5�o^R��V��{V��y��L^Zm�R�gٴO2qo7�)����N&�׫���h���Y1	t��#���deM8Xwl��y
܎M��4���_��c�ʎ��0�I���`����f��~�#C�X1��h�T��]HM��i!Zo�@��9uy�W���q��G`��:nk�߁C.�+rJ��V��"�9��3�{}�\WJ#]&c�n�}f�`)-8���?JOp�Q�.Ifƒ�Ƕ�!l��N��a�Q�CNMC���y��L6�� ꨅ[C�l��
��SrN)0��V!�6c�DS��t{	3̧�Q����\no ˜�]mI�})Μܴ^�}T�ט�7���$b�7\��΢�i
��V��er�����X�D-q���ǩz�`Q���U�m����I��۬ꎨ�(��Q��=��%y���QJN� �����iۮJ�
�V�(���/^m���Ʒ}]�OY�[zL�y���{�}��H���cM�#�����`�P>_�z����!e���%��n�TBϒpHx�F�L�}GH�y�a'5":"{�w�7��z,Kڟ��ʑn����1V�������O����S6����6�O��À���\�ii#ZX��~S+e��h[o<�a��Ѽ��<�?@v�ܔ��>ވRG1�q3lH��k��LRRB�T�]�����oX�����s+��Q���g����6���: _;ev[u�ɭ���G�YG�j�.w�3$�j��mD�s�RH�6�F���㡕���:���j,
$�*)��?��\�37�V�a�;%6>|��l����^�M9D�!Z������~�XR�$2CVa����̢�{��V�-������ʊF��ݠ�,�I029���8�^y�$8㚌�A������"�er�=�a��F���!������[d@42�K�uн��.�y����zw��sPOY�4s��qX���;��U�UD��M�;���LK�q�6�(!SX��I�M����%Tp�+�K/V)�pp��O��R`�"���E_\� ��|��V�:��o+]S�����`�^*3>S�`�"^_hSA���{:�ۼ���Y��1�N�1���u$��၀��Ԗ�5��^���fqkZ��9�-��M�ȑ�'/�np��I%-	�]��u�ko����H�!��:[B�+���H��f�c��y�ۛ�Q�(�j�l���4��6�g�%�![]OT�p��^v�^�,����Po�~��Y���_�tx�f�2�-{=t����2~I73X!.x��\�Ÿ���j�6 �:|�6�.�D��PW+�P)v�_!��
&��ez�{җ-�1֭Hm4�L�E�UzV���A������gw�����{�F*�F��igy�Dw��[�_����c#q��q$�����-St�����4�l���=st���y��րQ�YR�aM{�m�hJgX�y��pY1<y��t�e�zP`P��ڒ��T�h�*q��P�є}����@�}_.hF��-]-i�b��w��b����hKFE9�r`����!��un��@ڂ��V�QU�u�WYX����?�> ~���a�L��ե��D��&/�E�	��1W�ݗr^Za�3z�h�Q�,���A*N|���L�E�Kvv���"�����޽+�1�4����dV�%����4Z�� �D����d�X"~�w���<	��y9˩j�
�:�Ia������JuưL�:y��?��	����Y�<�6���쮶����Al��9�pJ.S���fp�{AYpʹ�M���Mh�q��E�tId��Mˎ��{�h�(�n���3�q���]��Ґ��`6�������@����:�pJ²`�Z�b�aƙ���dz���G==)<���2\-m�b����HI�E�vN9~j
�ǖ��Jm��A��7X�-	��V��w�[���`�cG�e	��9BXJ�\d��:#�ˎL��Nu��>��yhT�P[����������b#�F�enS�*L��E]}�� F��?�!6�_ |����9e
�P�?zXu�'�P�:Ih���K��)*,�Y����2�� �XY���&�@P!a���S3?~���KIc��
4V'�L�(�Ĝm���J�XHF9�W8f�8[G�q����c>4тOS��P�2e�h\俏k ҹ���v���t�m���}��}6�`��9&��;��jY$��/D�[(K��<0�B�*��31Ѫ�T�]Z��-v�nl�*���<A�z�ܢo	���JgksZ�/���ߛV���K�v���2�t���iW���g�
�J���hۉ�����;iJY�[}���@x��E:��W� )w�����e�
و$�.��L'�Y��e���wĒ��%�敨4ˣRJ�UU\`E�~�
>�1'rX���6����(�)�۲���Cכ�N�m�،�f��ۙ�9g���a�a&6ȁ��;<`��~	��B�w� ��-�~��!>n'��mƀ�׋X�-��h�O��Ug���@j�L���;�&o��g��?B���R���N�u15b9��)	�/
�VK� � ��9�dP�]��������i1�keK{d���<�k����/[��wh*]����A�_���ܠyL>�����[�? Wk�,��������TC��O���v��;G� �8L�c�����[/WL�1�i�]X��vP�sT�/Z���FV������_�ٶ��Hҵ�/)�����e7�<,e_f��z�Z��d��q�ɡQ��T4��7`�/Ӻ�ԚD����V0�,���l�W3DWa �����#l�8�>��f)�pV��9 ������v����#��&�d|���Ʉ)�.��z��v���s�X����+|߹�������-H��3�T
�F�b<nCde���Z}�^����a��M}@��g�&���-�H��Z$'=p2�E�o�*�#�����Յ�F,����u�gTa�Sp9��%���6�{���e]�#�6P5m�*r�ը����ɽE������ղv����Re�)�34�E^��`�z���)�O�̓��w�UI����%0{�eA��Ӿ
��4�I�_�//�=��������crڡ #�F
.n.��n3/���v��x*ēt�%Fa�U���km�C;��n#F��/k(�$	�#���b w\���^5::�&-t�y>�*Ҵ̴���-����Ôzo�]��n���|U���нo�>]��%��]�	Ӟ<�3yn��vf� �F��|H�����"U�6q�0�G8�}@ۤ�c�g����BQ\�[��I�o*���C�������� hB9�_�w��vAWy+�G�^���13�P�,�t���s� ݸ۲��~��>�BZ5ʚ�gO�� �caq���덷H�9&���^� P��u��u��OO�;A�Z�^[yh�-�� !��t!�:�l�@D�A��p��MƏ��|�(?U�b��*.�K㋻�y���� �S'��>C�-��v�4�����*b��Z�($�N�+�K7�w� R9����k��}�H6�j����P�4dI�3H���;�2ZNe"��R/�S�Ǎ��wZ��keB�Ԍ|9c�~���	���b)VG���o��ŻLo|$��8jTZ���8�	)<aE�s��F@���zY�F�N�u�[	��=���ɟ+����pzas�v��K�p1�`�n�y����%Ԋ:�?��3�Cu^����qλ�^g[�A4o�Zt��P�W�wK33��4�*���~��xD��!�Y���������cP�.طU��J��V�e�y�bG���-�v�R��֔5�>����s����ad��^�Iۛ2�����۷�@)Olr��V9f_)`���˫�E�]�~��P}~:�	�ꩶ����؀�?1-Pi�ٞ>��<��'A�N���s����Au1��W����l��[�s�ϒ��
�y~ހ��;31��#��Im� Y�IjW�s"+@�g4�S9+5����Tt������Ԙvu�D1j7�����,f���*?�@�T�JM�N��Rͭ�X�������2]��m��_��_���[8�ƽ}GO�$�y9��	��'vN�2���A=��)�w��H~7�Ʌ�����׵a��W'�5��q)D�i�� ���V�����o`���Q Lx,=I��Jb]�c0�.,�����]���D�\I!rHr�v3��H��JVW)�;�~���`�;;��� |`�D�KV}�k�*�pR�k��O�H���f!��S�߯�{N>��7O�]\�$߮b��5����4j�g#j����Eߝ{���	LQ���O���>l�PF�3�?��ʯ��R�3P�y%e����8eL�>�M���;2;�W�tZ:�{�D$ߚ(�Z���l�7��(Z>��5@l�]A��
,�I�5b�z7rX�W�AyM.��/%��R��p=����4u����jUQ5:1Zj�f8ˈL�:�$.�c��9�ȫPg�}H�{E"tcqC{X+���=A���^�E�JL���M��E�-n�U�
k����X�l��C,г	�9�3��:*���ld�օE6��F��J�������	�����ȕhi�Q�r���J��4�����` 8�ki��dߝ:�gLs�U{������w���t�@��&;����p�����G+���<�1��JNO�Z2W&Ȅ��~
C�w��Y�)BJ�Hs_�3� �u�)��v��M2���*��vN��/�v��ߋ.L�S$���+���t�[��o�M��A+K��ڄ��5�O�]����_�Ѥ��N<BT�����H��k&�N��b���Fi�L�=�г㹊%r,)���J��R�,	�I����4"s���\�2@|ϵ����\ A1����f�݉��e0�R<9�b�7QIq��$�*(Q�x��E�f�8qб4i�N�Yh4��c!y��� >�͊�����N���r爷�m�Y��w����^//I�����n�?���܎��?����y��D�}�Z��1��ϯ�"��d#>�W/�&d��9���2��3��`��-�d�p/�g1���fG����&��`���.����ʭ�(��3nڋ�{�T�@���c���$Pu

�}'�N�Oy3���N�9y"�r�!�?s��9J� �g����!&��������AO�p��e�
6
9IS[�df�WUe�ʵ�ߒ-|�]<�_O���&�hob��~����18\�M3�Ӗ�TUbG���)}�?0v�S}���z�C�ru�_Y֓�@�<�hR�U9[�Ȃ�!�I��@��TD��/f~Γ�ː��mگJ�	T�I�I�W�8��>T@O�s���l��c�B����r)��)LV���yRw~.�4B١�w���J�1��`��Sȏ���N�[�+?��;�j����-֘�m�g� �m�Lo9�פ��"$w��;|tωM�J�B��s�c�ӯ<��_���'����&V9N1�����^�1pM!d��?`�r��w^^>Qĺ3��4���G|^�ƶ�K6
�~"VZ�^ vʤ�>�Wۡ�p�$�C�u���-��I`�xe���੷ ��P3��w~t���r��ֻa����&�]%0�C�G��TX��\���;�;��"��р�3R�
���!�%� ��1�ML�S�����gS��<��Vz��`�ջ'E|�ɸmS3� 0�v�a�<ߙ�*���/bw���u������>'+|��~��WZ>�Yk�	����R 1���$dKu/��0� ���͏��2#E ��\�:u�xA��fh7*��IV�V��u��5�Y`��f��/o�P��;/������̳�F8<�� -n� D}$y�/�|`xS��������� XGmʠ~sc�,�y�dF�y�짬-P��Q	�}�"��lA�(���Sle�gt ��q��m��	���Q�`zg�F�?~� �X�_�k7��Pr��Q�*q��}2I�<ƥ���Q��� gc�;qU�{��8�O�K>9j�%�߽D���y9r�C�*�������M��`�QC��P��DI����9��L�N��7��U��$|�^�a��K�pO�Ay��zn���J�,n�}�PtJ�gGxyn�{�p�W֚��R���^���g5f�hˊB��}#ছG6�+a$���@P�ux�cmRK4�є.z�b{]�`�R�ӊ����M,�/(��+»J�+i�"�����U�VҖ�ijc5!A��u7=/{s���V^b�|,<zth�����������k�UN(�A��{�鯶9k�w���1�y����O-#G��5�'��kq��2�L&f���#�$�s��	������Ec�,՞� Z��6���a�B�Ck����P_.xA���j��������~B��?
"� @�� gl�[Pq��_�/F4띛!h���mH��*��Gv/.��H+�z��<� y^�e�r#s�15�h|铨Ҹ�����t��R�CG�'EB�w�8Q��
�L�1�R/�d�cЫ6�H����=g�����/���:Hw?蒟a�"��z3^�;��w�boମa�Q�	x�@�(���vɁ�4˥P�J����.S�]ݸ��|�`'�9��nQ+}���i�C�-"�xs�#b/�=�c��s�JKu��i�p��G�Ox����	�uM�o3�׶"���ޫ$��/q�73��h<3��]'��q@z��L׳��_W9.Fܥ2�J��~�X"�2�%4�ԊX�y��dnx���A�/cy�=Q����J_�ċY6��"���样�3���\�ՍG�T����8l@�j��;@�>���8�J#g<X���lo~����-�֨�����Aԏ��!
���>��Y���Ɂc�x��l9r��� H����v����>����	5���C)h���)4&��K�+�,�I��)B�B7���<F�7,�Ơ�0 � ����"C-x��w�	� �h�D%z�#cm��9�_��-Ur!��B�;��pRg_�i=�C�o/��I��i�@�s"!L��3G ���Z��X�jU�M�Ֆ�[Q$^�N�Y���w��J��B�G��I+(��X=ٔʦ��%@%��	G�o�<�A��_���{Y��:���=H��R��`��Oe� �=�\{�:���(���Ћ)
��՜f�w���̡�)��En�z��U_m���LK9�1m����o?YGK���8�O��.�|���r��ӵ��Lb�0�![�3O=,��y�m�2ɫ��$��b�OP̷��^�wv����pcF��[��RN@��T�3H��m��IL#s!7�!�K�s;l|�F���t�R�_0���8	��>b Р÷	GeM�7=�İk�qY�y{�$�_Hu�f��@���*�[F�d� ZA$�c�pk�,1K1���N���j��)�L�Z��aI?\?Ю���S�'Ӯ-)���m��,� �h'$�c��юsZB��-Ɍ���:
!V�p�|�޴����V�Oq�p�J��fb�f�16�Z=ir�42�ɒ�r��ݤ���X=������r�}~RK����D���"͐Ǜi���Dr��{{;��U4�e��uD*����=%��;�%N��nF-�����4l�'@�$���pZq �vB��l Ʉ�Da����-0e�������Nrh�M(�/
$�ӧ$�xH���s�1i�ؑ��=�~�U�)xS�u3{Жȋ�h����6\����l���W��J3�t2b����W'P�ֈ&z0�i�zs����Z������S���T���S����H���Oy�h��4�����~���i^M|����`Yi�;�j�w�:���u�(�<�����#IBuE+(�����r;��.Fʱ*��'d �p�c�y���4��͜H���?��7l��׼��xV*�[Z�'Ѽg�9Κ��j��L�Z���w��� Jz�(���9ovG	w�{��	�+"���0b��2O]�qJ��&����y������7/�#�/�B>��T�gm��x%�Q�y��S��;��ZK���>�K7#?!�i�4�+�]qwQǛ~`]>���8���8��;���*o�V9�o$�'�����ݹ.����Y\i�~E�U�H_����y�^�P3����O�@.�
nr�����<॥|;�����N��~�g�ߞ�4l��w�F�5�UL� k(�x8�q'�\��ص��������5��^E謻�)''�yt�g,X�d�.h����o~�~���Y���B4�e����\V���(r�m�$�.Ҍcb^��1��V���7�J��Gi&�΀C�iMkÉ5��h��(�x�h  �a�S��gZi�@iL��Jg�|�����D8�}�s�{A��a�;~�[�?�7�/��e'�.�TD����Q��/�N���I��-T*���:[r�tk���b7zR�P�r4j#�dn�g�K�%V5�y~�ۜu4���lB4��}"��f��e�9�R�>	<Q��aSX��:�$QWʹx�T'�Z�L�Aç�roX�Q�TF�c�������nH��	����b���D����f8��2<C����8Ű��a*�	�'*���v@ɻ!8�)g��v�'ΝQ+�*Q$���k+����(���)*J��?Yp#�8|}��qhW�^XP��>�R�3�
����(�X�[)��e���%'���bG�7�md���{�j\�C�6��W�