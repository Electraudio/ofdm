��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	�AVa4+طa?[�B�,��Dz�����Z�Wۡ�8ּ(���'���T��b�k�RΚr�Y��K�{�WY�VQ~��h~���u݈�[� �9����,����~,f��T�e��+�[���+ŀ��������9GL��n0	S͔L��k(�f����(�>7L����M¬ejܫ&�5'���R�^�����t�6��a��v���!���&ǄP�� ���=*~Ӆ�H���=���NI���H�`e�4ͥ��2����Q�g��.Qz�ffR#�EКMH��ہ�?� ������Ь!U�\�zW�#�qKH��3%��^�4��"��N}r]I��l`�GjH�]T��g���ڂ��~m��`���1��p�k�����^�G�ܨ�]�l;V��k��%/kAa��?0x0��nA�~hU2�Z��\4�u�*��8;w��E�6]�ǃ5��S���Zw4�c���>�ſ��S��7��Θ����>��OӀƿ��)O�� �0>�~�o�7��nF�
i �)],Q�����b�K��s�w�yR]�������l�i���<����>�/t ^�o������4&��Q�C�:_7��[��A}�[��4{��fV5w�A�u���`�s	pk �@ݏ�i1������=���M��8�,tL�`����]ؓ��w�n`,�?�P��R�b�U( H�+��|w�پ��LvM���b(�O������>`a�i���t�ڷ2��D���{)�eiQb;�ˆOP��v�:��Ы�l	�0���C�S�Z�e��`���_�k�n��N�ݤSG���Ux0�q$:�n`Ͷi# W>��*V�<e_�4��	����J�rEyB�u�9�H�m��h����� ��uZQ�bqՂzY��IAs�D1�z���u�Y(8���+%(�U:�Đ���\��g�DD'�/�k�4֛HP^et�g�#�;����������M���b�ӑe@�jl��4G����� ��9=��6�Ur*(�e�ƨ'��@T1+g�d~@so�~��$s�/wMߎ��df���?R8�b���QM6�IdXu/�E~y�I�d�YƲ*�ԑ}�����m�(҅��V�o/wzf�9{fktT�;1RCE��0��5�9�T��z˃�}o���B��Z�:�HŅ����F>I����I���:���o��9Ea]y����c��vK��sU�A������
�[z���2S/��D5%��\���ի;
��(�V�h�W�t�E5����N�0u�x�e0�&�S�q&�z5z��u�8fͷ�Y�<�w�����?��@˂�Y�����:�s�aCU��IH ������V�������+��l��H��(]�d��V�t�V�N�2�X��h!��%zj9�O��0�=��^�2�1���X��~_����{��n�$���m>?�x�Tz���O/��}SG~����{�0�P$"b�>y.{�$�	�4�Z+3�4U���	�]��>����S����"�Ю'�r&g���4�.��KZ����>�m�����+����A�	#A���1������-sNև☷����ZG`�5;>W�^��m�p]A�d� #J���LF	�	R�J2vʙ��n0Jp�`׆y����I��N"t����)Iy�f�&=Y��&�h��,���zj�y�;*�Y�:fo������S�<Ǆ��3]p oՋ�|G���0��3��k+�-���}Ⱦ� ��K󼇆��o�-ml��a���\2TW���ӳ���^ѿv����?�+�X/W$��Uk\�pW1)�R4.������~�T��+��Ɉ����S�م�Ze������5�����?�3�{���`�R����y��O�QW���fJN��9��(�5(�o��c`�]{�3	wz��ëh5�^��༧"�B5�,�����:dܞ����:�(!������ۥk�࿠#�F�^���^w0`����M��B�3&�磨oQgq�使��,d�l��o�ׂ�}�OC{��fJĚ�;��J����ؿ�Ev�ڿ�5�G�'��a���%aߠq@���6Vh�����:�i	Hp����96D)��T��շv⑸+�U�R\�g�u}e}��Ul]��3S���S�*2͑�lUe�?bW�ML��%��bL��]Ls�MK���f�H�jݐB��@@=:�S��`�kc�~Ĥ�P^|p�0�b��H���Yٵ�x�OSv�5������I�$G���2}�	��0�s~��i���!����>�j��e	0�f����C�r�~DD�o�bG��1�^���O� �D�z��*��l0ޱ�!xg�Oň��~�+d����H[zAɆ'���Q+�����4��ﶪ�R��#K9V�#���5]�٤�T�6E-b7��;�m�|d�6��E�n��w��XͿ"!�a�tj�ѓ�F��&�p��vc��ș�Y���i�,�F.FQ�,Ĝ�||#������{:����𾫁T�]�3ԕ}��]�Q���x�*7����7i���0u�����=��T��29�G���F���%<��Ó�.��YN$�ux?n��Ի��xI�u�9��_����ܻi��Ao��W�[��A�U��Z��G�l���:��M��VIa�A%4��ណ�ܪ��v�CE����P���Mѻ�� 0�A�?�(�\23 n�(�#�Ŀ�y��t����=�����fw��'�FS,	�`-R��b��q^ٕ&P��8���`����8��@�s�I���З�ٰUMs-�#VI_���r�%7��PK���׼�TU� �"���ɉ��]����S��>?����t7�k8��N3HL�z�>��ϰ�-�$G(O+��s�g�[<xm�q��Z"Ӣ��ٌГ�Z��n[�����4��N�%-���İʝ�� V؁�~h���}n�x��ׄ�ϳv��ҽwi�T��1�/��yj���_%�{�!�Xy��̋���0x�,���q�	�õ��z��u6?ͦ5��z�[2.�
a�-Y��e���~����լ��[��`�'��`�:� p��]�"�����.:9�z헮N��<�q��j����jI�8^G���֭P�c�g�u2�ɕړe�: �����|�V�P�y
m�"i�� 8�����I�W��.�q��V"���s�su�?{����]��w�һh�q������5t ��x5Ps�tm�x��<G�t�^�iȜ��?G�AH>m��Ǐ��`?��"/�j� ���m��O߂a�׋�ƍ$A��^�aѽ�}��6�A5j�%�{ϟ���+Snmi���Uz���B��vf�%T>}�K�O�&�;�}���`;D�l���}���S�Q���л$�PYx�1��h=�����6=]A|E� ����Dc��CBC���-���Ǫ�X�:�����7��u��Snq����+�:q�G�{آO`�t,f�����ˍΉ]Rrr~%C�z��<�=�ӟ0 ����}��\t���3��/����:@\�Tx-��:�n�?31JF?��%����Y>rX4��<����`�-�o2E[�\����h��Ak�i�ii�Q�[O [ܗZ������D����{�;���D�k)��9e	e?ǻ&��0��ǖ�-t+��U�QU ��.�9��7.��-^���6�b�z/�8���*A4�x����O��l�M|��ׁv,x�{ڏ�Ė�˿�e&>*Z�
���p��Z�$��`�����Ob�*���i"�YW� "�%�	�fB�@8���k-6��W�m��z�΀�i�3����ʮhB1�Ѭ��X'�	o.!�19nʇ����ߥ�@bK(���K�D��9���	��F�#JR!p���@�?Σ�����ܝ�vs6La�z�r��2���ndI�+�F�HvC
�S W�$yڃU�|��2e*y���ύ � (F���o��v�5��4��G"�B<�m�ʆ\�j�Si���K��"0Ϙ�l�s�c���eay=�]�")��XɌ����0����Ϫ��X�}Cp���J�R��}y��͟�P�h����Zjh�#�K��ʡt�P���w�2�wu&Y��� m\8B@1Q�'�"�n�&PDЦtˣ�q������$t��Z��RT�;�yވBf+��5̙�LujA��\~h~Q-�r}�+Zi��m��^?����e[�߶
n��J e�;f]폫����o��p:G��6f'Ĕk��RV�,O�T�G�HsGk���G�j�9��ИgOo�'9����r�n=e��O������eR/�=ڪ�KZ���M$��� Jx��?�'+�q�6���n?���*mr���U��#����}T�S�M$D���
��W�U��������s���5�5B@�OAf��i�����\�Bp��n`�,���<�~Kt��h�qL;|Pmc�R��o�M���U�;�d�f�\H��٣Jst���6���Z@z$�g�:�p�,�����|S��@l͟�P�.�Be���At��lD� ��� 1���:Vf�͟�B�^{�Im��;�lv�M����E���ܲ�=�>����	���4��*���t�A�=xP�.L$��
J:�ã�I���S~h�-�������� S<�,a���W��ù��,X0C��_K������#L��ՙ��.O���qV{i�.Y*�:���+����gF�x~��{��8��@����]���7LĴ�f�����Cv��:�~0uB	1��}�m���.X��F����=�-�����L)f�����������.1�
I%�2. �ݵ�����������e##2<J0�9Ȝ�UUT�(��/)�m��^^�X�3ϙ��9���}kWK1@|���]���'Z:)D���
��9X^Ӥ�r�gP�R���|\w�gbk���0�'�^��ҁ�!���
�=-��!�a�\W̑�
�hx��� n��#�YK��@r��:S,�PH�?�Q���m��<��j�{0c1��������W�>���bTOp�!LƿĻw#s��
��r<P =�U*���"�fcv�HLݱ6��ܘ�{C�1f�i��>(��~Q|tF��Z���'t��}���h��H�
�0m�����4�N�f�'^��}�^1�T�o^|�p���D3]ʾ����Õg4,�%��%|�xW��%��4��R!�Hn䵝�
!pH�.�Ze{O���C?� 0Yۤ�4�#���R�>a_s�=ב��$�#�=�96�i��>�~)uᠤ�H(z�+m�X$J��l�	��TE���)�[�(&���,�W����zs�j�� �B�M�TX��>A=0��I,`մ<�J���ߵLj�̯���L�� �^� Y�m��;݀�L��G����ٵ�p}+�G�r�>��/�,�P<A&���t9�5v��_����xd���)����D�f��+��&a:#�R��aQ��x��K݇2��1��� ��Z��^-V�2ٗd D��-G�>�cDh�p�3���x�4ESa�.����CL�*�w��ը��N0�F��=���1F��̆��5��$C"���o�К	��EF������������w��Miͣ8B-�{����%���u_F��c��TJ/����� (�QV����&����Z6L�ؒ@D|�6p�	I~ƪ�F�� ���,��D��;[���7�׏2��P(9�����U+k+�/�sn��S�w�ܼM؀c�ɾ�`|ݐ)�u�S�����rx�Ș�����q}��p*D�y�3�qt��_ʕ��qB�t'*�
�{Ґ��P��g��+��!v��w���տ��mZ�>�<rh�0��<y�l?��/2&	��G��RuA#W�1����:�1J�slQ�
�?���s 2�ur���MF[<�`�ܻ��0Y�{�û�J[2;E��%|XX�T�c��3i� <���$��+�4��R����$�[��s~�D͞��9z���넳��PV ܑ��1rk��k:�B[�3�uU�p�P��I��E�b�f��0$/�dE�ed��R%$��ƫb݇O�'(PX庴�Ic�MSz���J��O��l��AO2Ӫ#͚+*,�ѧ�aը+k��u��g��G�v���H^<s�+�U�Pu��	G�Ni=�`�>���.���5N���D��_hxjJ�R�[`�p5ů�����@�N�*Sީ������h&B<�4�JҙJ�&�m'������Ů��W
W� ��WxӞܷ5������
����Z�Ȅ\��9*����
���G��'�8hH�Z;)�aGK��}�[M���׆��Y+?y��PA��
��i!j��(oՃ��9�g�6/r��jC�O~�X@U�8o��z,D�<����Ј����]�U�Ot�ҟ�j�3b��*�Oo�u ��������zo���˭8�'��︾O�)l�.�-�T,�rS��S(�ڑB5�ێ����zCN5Ŝ"�u���&.G���&V���9��Їs��a�����������N֎a�C�����߾oj)Pm��(r���C�����ա��mi�7�}�p��`�v>34�%�2�_���g�4b,Rad�����mۘք���]���ޠag�4��RU�j���}�v�-�f���X�����Ӌ�f��}��cIP�W��f,<��.0rI�n��>�Jf������?��Z=~rRHgb��aJ�ދ1�t횪��&�pwާ�yo����,�[&9� ������tS����F��c�{ʘn9�X���O7:�=���YlΤY���r��GW�3��'�ÊMo��
�Ҟn� ��	�\��'�j+j4�R�o��*���*�x^����cמ����}[jv�:�a�Y4��-ː��Z�|�l��4�wwb􏦵Ac�o��5�0�4c���
�҇�p�wh�`#_Ѻ�� ���R/Hg?��y�0�����к�7iфW#���E
�w1� ��"���h�Z�Wc�f���0�PܹJgu�#a5�i�D�U�m�X�t:���EC=;�<���B��FOX�k:����٤��^����>���+��1"�Ԣ� ��5�tv9;��ƞ§ʺ���x�Xht��^��{k	��&Ϯr��-��z�?��Ψ������.�=c������ԁ}��0e��0�]<��kf����=�cU�8��Na��ers�������t�4��m^�ą��C�Ń;��3���h�y;G)�5�(}$��ڢ($���Fj+��t�M�aFU��Za4�m� ��)�a����X��)hn=��)���]����t����A/{v���	��G_{�N��u��f6�>�V����ԋ���6tV�-����D�7�0�E������FP�4��� 2Ԙ�Hl�f�~�G��xR��B���(ؕ�ɓ��kZN�(Eb��p�`�E��#�[nG>�'�>�p
�[LQ�$:ၫ{ۈ&43�c5RQs{|����ʤT���L
y�I�IӾ�2<}��!/h'��<������������O�$�R�؁.oK�����8��}{Y|�{�����>�k)����Q�����\)O�PMSNt���O�S���ϙ�2��0��A��TsO���Ǒ��"����,^>�DW�
��%.�*�i���oDc�m,�y87IU t��u2V⮒��fK5Z�H�i�~�<^LO�7r��~��o��J�F�H?1��S"�h��(9�-����4;dU�#��G
 �����)�;�ox���)�Z*]���AA�#(�	!�i�-���z�m 6+��+� e��m�"�0TUd��&����R/�F��{<�c�I6i���;��d�T���s=�V��Y�q��mx@�b͋?�zr�����;�����=O�"Ak��'�G��{��I��v5/���+l-��6�<hl�߷���Oסҝ�k&��W����A e������⟿n��|�Z�p������8t�;%��[U��X,xM9���x�G�f�Dz��xP�u�ϬP��Un��ԩn�����6�M{��8��)��R������g��(�w:���ݨ��M���err������͠�bUh�:���Y��Z@��v�����3�����?�2�Q�5U��T���j3S��?G&�d'n;'��S���	�����zJ���� Z�,�f��_���nd(J�����.�j�b�(;%���yI�.�9tx�G�9����S�ǰF� ��6%Pv7.6vb�l��CM=e��2w�dK'���(#<���n�G��rJ&^ȯ������ľCHR�Ů�]�;J�g��&~+nO�Z�T�Z����"������jJ�[�V�6����C(ˌ�+V���%��p9*�&u��E:�+ӆ�B7��_����-t)>P��e���F'��:ݥM�������x��a�!O�e�e�;ED��:{)iՀ�Ժ�#M}(�Ї+پ�ǽ���Q�����;nn2��ne��r>��#��޴J�SЄ�Jְ�jQsHOpy�AԹ�Q�v�0 �/A��`���k�b	Z��f'������瞈e�w� �.��r�A`�v��ޭ�mX&��ފ�LA�4*W�g�m���Xe�	]���_�@b�0v�e�l*4�g�X�՝I��^"v\KM�[%��(��o6a+�²��-=�b�$�	����=!O�IU��2Ϲ��$�u7���L��ɰ�L�	+R��G�3���Q�og��M����h�2������S�=�h;z/�R	�l�x6���1o@Z��4BU���T�m�lbF�9g��~j��<	�n�����xoA�/Q��.���,XBX{�j"�={7��9��N�~��U���O;�^%��9����Q�	ً��ԌG�4���9�
�@���y\Հ�A��>|K$�|E�$Gqד]#T.Ҋ�C��$u�	��wS�N<�^����׏뢇4���Tw17��.PB��9	���!���cJ���e���{�B�)#ګ6�u��CnV���iJ{�Y)^E�S��ݳD���2ߒ\Z���ܑ� �B�t����`��g�`���~��J��v�}��wk�}9�]qnĈ�Ѧ��x9Sd������0�Y7�lc�b��Ya���%�b�1(�t[d�k��,�_w�+��	1�m���ۏ� aPh����=q5$��������ךĆ(�BM<�ܫB@��ƺ]���' Kw{@����5`@w(��X���.=+x�dn���s���77�u%�d߃4ak<k�]�P�����\_kci�	����+r��VW��k����{LO�>s�?�|��S� U*4Yp�B��7 ���� v�/B��K�+�bF9�m�끤��:�Ra,���� ������X-��᭏iI-�J�pW<Kwe�D��D���c���=�G�O1��E��� �"�*�t���� a�Ҍ�C<=AXaE��4���nm"�(��������ҷ���B-���+SyJa���|�5fh:�|ZU�[�j�4��sٺ�ϒ�h�QŦ�t?w�R�rM6��{�d���8鳪 �r4l��]*\��K�4a:�(�h/G��X�C[����Ve�cMw���$��c������ֈ�"f&2x��Аl����}1uD��x�wyy�[�n֡d}�����x�����͇�2q�D5�����V��U#�d���Y��X����bK��\{H�=��O.��Fd�;F����;���ﷁ޲��a� #;�� �a6+��En��w�v��?k*�]69��������U��G��xV��f�UhGURQ;��kO��q��?��O����M((�B~�,����Ҟ����{���o�Pm�B=��iq�˺2�B�-���c��,�Bu�V�9nd�}*m�<nF��HH�h�Ao=V'��8��A�3�@�������<�SN4n�.�7�L�|����@��2��d�L�В 1d<p�hI��e�� }&�����ub�׌�RxM=e0��9j��痬Ɓ��I�8���N�V�G�\`7*��9�~>w��,Sfp�g5�,��4�mǉ�75YR��6���g�����cw���q#`��<�[?&D_;,3LI��/���AS�3�\Ņ(ܸ� �Qf�B��#J�O�����Dض��Q)�R�`�<�Fp,���ɦ
�/�S�*���(%��R@��2F��{����f5��e���?Z�Q�����?�wԛ�BBx�`��06j����=��I�#�fm��a��_/0Uټك���)3���gh��}%��M*S�}�]҈^Y4fZD�n���RLL�]NW�.#⢋�Q�� �N�ˆ�����[�Hpi{���2�>>�G���x��o��9L��L���ʹA��B���p�I�<Pv(B�B�5���Aq���z�ІǗV]b�P=N�<��o��kݴ��6�� "Q�J3�7�EKw�j�x��_���ի |�6�%�����#I�`aP�牋S��oA0oM���wz��qJ�Y��	S>�����*�����o��0�!���y��/��n�VH��WD/�W1�������m�tķ�r�W�"tG��3�_��לyƏ<F~��r�+Z�҄�Ԕ�W��Iy��##V� ��Xe�Iq�_�]�ki#膝-A�5�n#8_x	4T��Ҕtt�3����=X&��E��}�05φ�IY)J�J���� 2��N�:�t���B�R	x�I9���?^��`���" ,'��;?�%�k\�W�Í�N�М��Lg{i�~�\�M^�[;�\��{O�w
���N�&@���-Ū�Sȍ'6�Bį٩D��#X���w�U`�>�q@T1�i���u�O_/A�R"u�{r[��S�>l��8ӈ��rA,�%Q�`�4Rގ�k�˕+�&č����}�l�Qv���M˜R�	˽����$*Ĭ�X�m,�P���KL/��+�E`��7]�w�p���K��4|�g�fX�;!HSP<�\�t�<hKQ���}&��Uǖ�j����c�J�D��v$$ed5��o��g��)1>����HS3�SoU�#Mv �j~�Λ�V�s�+U~F��������*n�U�A���v���/�s�3�&hGϯ�.>D�p<f�
"���nF��$<3s���+[�@ŚdL.����8��Ag|Dmb~���q�Oh��1^����7����h�2���o7��/ilÈq~��=� >�4���m�3��'��IR �b�,3���#�ޕ3�E_]�H҃Y�\��W!���Wa~ +�~m��7-�Dǘm��s�]�,�Eƥ��'��<'���DG�
��F��i,���"|.������
{"�n�*q6pft�I9��o[bn��nӒ��poB�}z�n"�j���yBk�f�k� }��?��1�I��=�p{i��``�֮�|�X��A�P��3�����l&�9��5���(y�R��`[Kg>D��|#��rr��eX�:�]ǑxVω�0�s_w!:��WR�����]�mfѻ��Ϟ�֯7��Z�+��|��A-5�����ð�D�,��Є�q�����*��T%=�<.=q ��kW����7dq������5�,����*,�ZW�@H;~64ey���d����h��a�>�&�o:�u=8���1�vX��_�>nÈ//��G&�¬l����R��eߙ#9���6F���g���
�X�g0�b�?��<��}>�sm7�d(WV̢T���k=�݌�c�����o_Irll���q�� c<8�a��2_rG-�qo�Th�Qb]��^%�=0�"�����Q��V�M�s{C�@^�t�}^��:� N��Uތ,��On��+��{uR>>^���n� �VϿ(�S���Z��67_���O�S�H4��F��H�V�9lPD�^�U�QJ� ��SB)�V���`�!��=��b�o����Q�H��/�?�e9ym���0}Ba=��}^4�ȼ(�d�q1��|Ի0��Lx�S��1��8j����yn��+j��9��͹���5��C5#Ym�?q�p��C�N��������5�FR
�R���(D����Z�f)�SW� �Z�piW�3�H�{�ك1֬Xf�8��қ��[��p��F�N�W��^l��H�j���;�^r����n���쌷�RHᏉ��C�q���כ�0�a$��:w����s#����3���H�^*�״O����B��T�]���\�"В�A�"��� �*����ץJ}�x�}�D��D�]8S��Bm���9�������Q�:��d��ǽ��;b4�7l��X�kg�Ѫo����{�+���z ]	S�_P�&y!�1�de���1�`�b�L�
�
N�%���^�'��;�pDN}ʦi����̘���(��;�P�0�?���fP�\WVQ�㧃��:����c��]ylǚC���"��q�o���DfD�IC��iJ({���0eE�I�\8�K��P�M��r���{�{Ý��A����ȩ�é/��mm�	0���a�<�����M�gJ9��|M�!F�q!1O�k�A���A�<P���C�����.R�+<ʏ���A�_1�&��-<!.O&��6;T�
�ܯ���k�Y�v.Ԑ�d�:�+ic�����6wa��9{+��j��$���xQ�Ơ%�I�#�D���ҁ]1��{D6d�B.jL���qS�Rٙ�\���"m��[3��W�O���4G.㵷��Fd�n�.����0ٛ�G����s�3	ψ��0��{c�ܘ������8o�����vC-�'�g,�-G��cK��R8b]A5Ԙ��h f�S�l�Q%z3F�;A���xG�68�g�W�4�D�o쇅�PE�ӻ<�項6��r^�*p�x��O��OE��n�.h1Ww�TUk�\���K�X��.M���x��o�C&.���b��++r�6�LS�h��nEW;V�����O��k�rtl�XQ�_B�&'Tqtc�k�K�<���Ղd�6@�HZ�H*#����*���_�7}y"���n\����M��UG{��芀M!��P�c#ct3��,e�$�P����Ɍډ3Ǝ����d��f�f6[���i"Vv�d�x��G��@bAbX^#��8~wb�@�����c�(�Y0�DЌ�19��[���^�h�;}�-*�1f%�zzd�B�Zt���T����ރ���X	6��"��֪	{m��W��n�� a�./۶@\D��R�?�1�.*�ʬ7?BD�D}��ӓ�֡�5��aZ�Hd��T=kd3T,�r	�h�"H!�/0�	���q
��[�{[`��� #>Մ�����'������y$��SH;XH쫷NiM{��y�����x����;�-�T
���O��tg&Zq	�Sn�~B$���#���C����*v*z-M��;��il����e)R���V�z�.n �NM�ˀyo����qkjN����0�&w�I�(�����o�;�������&��u�&�iQ7ůh��"W&��آϝ�)��O�����]v�j7���)��z�}�HT�x%f2Z�-��@?ʩ�!u�SF?��9��t������"Dx�q{�����'�M�S��a)Z�v�� �_���{CϮ�vS�� ?44@�a7��4y���/�q�J���,D��&!V���~�A��~��\	(�8,�;�bD#�{��1��I��P�.��U�=�����ފ��� �x¿��3�ճ�g�Q}�?���&G����g���y�	(s{�\�_�ܖ.y�Y�3���GfPF��� 0�<�⍀&u������/g%G����W�T��j�C`	=�yGN�1�W����/��NQ˱�v�0�k�'�2]�?V����6YM�(;��=�f�$�dEMZ�U�?��J����D)?ǐ.�m��_'c�o�<O���륩AXӓ5���Dц��Sݳ���w��U��,���1��J5�����@�3���y�lÓ�g<ܻ6h���=�K4�R��o� J^]䳈6�h�����y��KH:0��5�u��j9��������Y\Kk?�w���k�@m�j��F����'xF,��m�0�e敛 ����m��ؚ*m��x��R��R�F"�"�!Ag�����K4_���� Բ�_g/Y�Mu#mG/0iڌ�â�ط��.�Z90�h���H҂���^�>�u�3�����rk�F��F�������9�T�I�Ǻ"�n����������:d6���_8������ �J5k�R^��UN�)0��R��1�6R �5ǛcYFR�S�{Dm�}!�_AH��i�~e�H��u_N����_��4L*N�[*a���Mk�f
�[�48l��\��j/dV�����{Y��U���s�y��2�N���ڮ{��E������̂���y�uf����E���0�-&�H�V������7�����M��d���lVa_��l>����.���)��Ɨ��:A>�y��L����͑�9H�w���\q�w���*v�H�*�Vk����X�rΕ~��6q�d 1}d�P�p��8��R�S��-�`��-V	��	�V!�g��1���V[�(7����ðD_�V��˻	6�N�q�h��^G8�&6��ǹ�6�'�L`�0*���� �;��nC�T+�5j5�C��� Lyqo�#z�Q՘�JM�^���X�p�{Gs�����?h^�Z����D��9�L����~�t��ݟr��Hi|ۼO۞|{������eŪ�7
!���3a?�����a�D�I�{������٧9�� ���T;T]EY�ԗ[g��:��/3W���/{Ot�8�_���R\��ͷ������x"�wL�d�ss�� ^@���z֞�#?��{��T�D�@N>�	�N��w&?�N�ۈ�6�7f�����'�̜ˢ��j6�F=*��8]�ү\���
/����e�I"Q �3�h?�|��*�g��Mrʞ���'0}<c��ܐ�Ϗ����ghKY9Jjm�ڻ;샩RĊ�P�U���-�ڞN�L��d>��I�-7�p��d�n��̉��+����G�*��%p�v��#���_���J�PR&ދy�cH��|L���#��9��m������hal�������"�^���^i\C����R�,6Y�����D�ѽ�Ȍ�Υ¬0B�?��>���&p�4}�@���ُI'��2��������i>�q��*�`>K';=�i<)�âm�ْ멲�p��_^��D^<��=uLyG��M��G<T����K�P�49��|�%� ���Ck����^7��pi�̚*����>q�&�^
}/�i�r�����-V��L�2mU��ZzUz�QY�戀���9-6u�D!��rY$o�/n#����kl�/o�4�S���I�<u�V�|�� Hi`6�� ��t
<��.�yx�.غm�>��4-�j���R�iD���u��DW��KXd���i��bK�1'��ɏ�-�������yQU	Զ����/���g�]�r��_i���?o��ʛ��v��K[�| tE�7���Mt��X��/�&��͢抯1�����bU�iP�g�:q Fp�NZx6R?������Sʂ��ڌ;���F��������>n0�~i���g��R�;W��eJ`6�J�F�%���iCL��O����_��*����b���+旈B��9�+�J��2�vh�^��@�ء�]"���!aE��׍P(x�8>R��]j؆ ö��od]���h����΋�C�����F)٨o0'��Lbj���")��j�(��oѿ��ˍ�ê�L1��Z���^�G�n�qm����H�>W勤�����@��l����F��Y����
�N?�C$]%�.�����C�qji�GfH���� E-h4U�����e�y����BM;!�n�?���F�I�t��,EPŅ�q@&r��Z����އ��n���9�\�`���#���TK;�. v5E�O�r��i���,sn8�
4»f
�cUА�C���������G�����K�^� ��ҘB�x�R]ߠP�����ny������>��:f�k��?|���g�P�;�~������{,+â�L0�R4b���CA�9�L�1��^d��d�9?�Z�c�d�I��Z�ۂ4�r��:KچP��X�/��#Ѹ�~�rR��bZ����l!e�]��t�â!G���V���
i����XPQ}q��幎�i�34IX�,�ͪ�����A�?���8d;����uL�GP7�(۱��L��Hqj���ᲃ�����ǂ�d�#�$�rpvt��:�ܰ������9"��K
o0a���@g����<_��׽s��9񣅶
,Ű�/��8Pz�3�]43�Ҡ5�,]}XU^ô��t_��^��������1m�=N�m����-���W�Na�-�� (rLPL̋�a����
�7���d����O^��Y�']Qo�l��H���=�iƍԠ7օ�_�Gc��KY�;cNzD�ϼH3�y������7���4E�-�06,E���t�3��@���ͧ���ju���w���a���٫�fK׫O%f�(��1�Y_Q%�^�����6�R�}U��`̕��o�B�����\ ��]��H(���O�AL�cH=j_�Qw\6Cߗ=H�Q����R���o���	�kc�l�
��E��B�q}�I�2��l�'C<�[�=T����L~$ݺ���[i]��^�e�G��q�3���o�a����a��E��Ʉ����TT{#�0h��<��)s;0�x!��@F�&�����-��U��7L���Z�3=���ixI}A9qU����*��ϥ���qE�%����pe�;ZF#�K{s'��Q35-�Ϙ�|��D���0�8�u�nQ�ZҌ����%:K�rX���wk f���w�,���J?\�e� W�G���I�l�-v�E��B�z��N�(a��Z���T� ��
�y,�E�5$J}��{�V'�|({Q�$��t���_>j��$��6^��,����OZ�����V�d��N��/�d��ہ�N8�_B?�R�wB���0�,_r��
;û�yZK%
��	�-Z�(���t)�t=q����c�m�9T���ED�b�y��1�;�{�A��*�����!+�v_��^�ƜF�����'=��S�W��Z����s�hL����7pN�r�a�����h�	���}��Ƿ'��opF�y���|���ϡw87�S� ��K|�N�e_�*��9N��:����`}���Pj�c�� gPpcTLH֖�ԹA
�"]�b�K� ��DG�F�%��7*1%��8�B��Ȇ@u(�L�Z��r0�H L^u�O�5	�#���=pvjԣylw����L�_�P�'��ޑ�4&��t�m�3|��t��u�Q;c~	��B��Ro�3��5�S����Nq"��������Ѹ<Tw�dz|r�3q{��կ��bkQ��,݊#Jp�bz�֯.O�m.��Щ�C�Fy�!7d��l����2I�<�������A� ��p>rys�ua�μW��ڠ<5�j��Wh�Φl�����a�~OR`0Ȑ�\�?P�	��K]p�ڎS���Fŭ��D���-�ק�7�����ó���FC����x5��<�+����xj�W�Ч�so/GS��N;�>�y�Qy�h��ґ𷤳�p�����a�uc� u���	�	`���)���Ҋ��!���Ka �So|/O���QrdB��=��7r��j��ݓ�"R�ܼ^׌3Jke�XU]Z�C�������8[-�����������<�x����$Y@��Y�[������)H]\�����<Kiie�GD{ِ�@�Pa��/}8M��%�����Oe��d`i��l6 �2p(���(��3�$�?�bKc�_��}������2`��5������AG�5�/99����Zao!WF3LR�t#������k4�#�Z�*D��J ��la?�N �D�� >��A�>�P����>�Z�{"��U߫����]��A��W�ܨd=�"�b�����,��:Jv̓�QOf��h�:f G�)̼v!��u���������DqP@���E@��HmQ���\�g�D*�
��>
�c87�Ը�K �aI;���k�'L�C����<�3w.P��:rU\���gh�P���C�S�C��磂X��oN1	�2-m�x��w>�h�K-D�X)f���˥�Lh�fщ�r&W�Å����pډ�A�U������i�t>�g��ԁ��y�!�X�:�J����!s[�f>#�ܰ�Ò<�<&����T����M������[��<�*dbpt�
:�_���rLP��u��3 ͹��L3��]z�@��(�)V<�Di�v��RΆ���׸~}:�x;,/E4��z�����g�ˌ�ժz�����BP��b����궥DǸ�)���Q}�\�N�n���Qx/��4����\~��湨��W�@��N#���0�}���s�s���h�0�?��)l��O� #d��J�L�s���)�����L�^k��d��>�g-q������3& װ�Z�s������	7�q�mY���9�{�7���6����os�{;P��t�<}`O^00��06@(��.�x�kK��2��?�|�zEV9�9d��Lѻ��}Պx~I/gx���B�S���5�{�Ch7MSvǎY�;Q�Q0��D%���X��3�+V�u������/1�6ܶ{w�yc,䕲i���Y�b{;���n8���A?�A��a��MQe�A$����yOO�FzL����]em��:.���}q�h���w��.⽱Үۧ�E����Wpe����}���ؕ���!�E�pTE�����;�I��D�աK*}=�4����QY"e�A6�t[�./b�m�\Ϲ�2��[�H�6�Z�>��d�}�sB6>u�H6�ٵ�d��p����y�!N+,�֬�E�K��6
�2~|؛����3#_�a-�}䦤��+����r�V!�y���\A���A�-dUBa����T��%^&�>5�lO �r*�Q�T��sU�)v�|B�7	�ʴ�J��gJW`)}9g�6��"��.�vW��SĨ�͢�*m�0�dA"���I�R	�G�)=��$�"9�[�YqA����̝nʸ�_��62��B��@è|Zl��{Pښ`+��1�蹗T��wi��ih�0�����W޶�{��Pp�w�B�?�:I��#X��8{[X�+.(�C��{�kK����;��*���/���Hni�%c��+���_��o���B�'Z�N��{<e������6ja��]���m.�i�����B��C:��r�>Q2���3S�`�K���_3m�|��er�=��M �H�������l��Dx�7?�x�!�K�G]ݑ�R����?�RT�	)۴p�����,�ߔ�s��Ic�?<��}G`Ȑ_�Jm*���#/��r~Ϸ.�901����g�[K��aW�'������pӫ�����	7�[i��ZN���� �����Y����cQ��JIY�_��7��3�l�<$V ����&V��%�ȗ��V��j��WQ3�C��VW$� �Vf{5�%�A�l���������E�a�'g�9�7-����N�����W-z�S��T��&�亗���_3=gn�����������C�M�����	��-1�\-��c����#��~3�i���b�,��O�}S�B��:T>�l~V�-�}�~m�M*�qA��m�K�K֐�A�x�w�,��JA_V�,DY�=M��}�[ÞM�U�,T:�v���;
���j�����X�uC�Fj���_I^��]���ʒ�mJr�M�m�41�ei'��0�?����Ȑn*� CR�W�u���J~'�oq�����ұ������ m�1�"$V�i#�=�[d^��u`J;O�;�my�\��ֽ{`]�9	���~[��9��9
�M|��U�CUi���(W�C�����W��i\m�
��f�PG����K�� Z�,S�Hi�>���=�qnWz�U�ƵF\	�b4	.��O�����Z�G��)�?�(�H�K#s+ڔ�X_�f������w��8�i~\�0߯�� =�~� �L��6�$��L����qh1���->��$��)p��u`�B3I+�bAC�H&ZP�g*:�_��܎B?>b�L9�l2�u:�:-�x�.�y3狦��g�H�a	��G�9�̈X(�a�܎�䏥�mkmF�;(t���0���;ER�f~��St�Z�`�T).��Ӗ|?��Va���*;����yȋK�a�&����#�#>K�YG����D�O$����	X������3s��,��g!�o}�ǰ%�6?>h��T���8�ś��O	m��!����O4�
Xt%�d6a6?/a�I�'���]��\c�Я�`>�B;��2�ɇ5�����Mϙc��0H!�c�KO��신�^�����x���;�(}������:��W�S��1�=���*`��;F9���l�-6�"����N����j�>1�AK'� f7�Z�O{��8�vk����	;B����ntls��U�?�!���e�d� ���w��vB }����}Ij�9�����ǯ�[����	5���Bu��;��rM�N�]H9�j8����/��՛ݷ�:��٢����L3�H��
?U��I���,��*! Ü�9�szxe�����R:4x]JU�7��C���w��/�Z�.�"YT�I' �Q��}$g���V_yY~� '$�W��c%b+ 0��,O��<�y��-�X��@��:D��GE�@+�T.��X7cmC���@䐄n(���'�O�v��퇁W?:X��>V^�*fs}�G��jT˽�C$�R>C�|+�/&މg~�D.�K�b��5
��[.���k�4��Q3Ⱦ�ܭ�0�Rru��w�H��������s�gN������jy4$\ sRE1Ư��;k��F��HObo�%q�M&]ޔs��J]�ëgF 6Mg������A���Q�� �O�����MQ����V �J%�I.���9��=�]
OJ.���WL'_�������h5�4� �5��J�}	�����.��;@��)8t��n�Z.��r$C���ٷ&|-."�?	�d-��Lg�OYs��L�^A�šHT>)��u�O��`c�-Q_�z`����Y�W����y�7L4�l(,�Dz�
�EDa��CB�t���Ғ�h�i ��l�8��2A�`+���y4e��~d^�dTf�+?T�V$H���ݰh����L��6a/:X�Z�s��@�2I��<fa�n���P_�I6�c����O����, o��B�I�.y�]~����,5[W��B�"-<_��[z(j�KhA�w`|V����f1B;�tjU~[�Fς��c��G�������w -?���"x ��4h��[wW=�t@�+8(����v-��=�i��.�<��9$�c8�С�4����w<��7ׇ"ﭿ%��?{�ӂOP_^�� e%
�:��w�G����ZD��m��� � 8Xs̞\ޞ�z��/�T�˻Ņ��Ć���e�@<m2(����ie��
��N�k���
�e6��
�!!����C
���0��ڕ+ޕp�Q�v�(��:@*U�x#���^��9�˟8�Ƚ\�4�К��}W�ӱbn��X�9X�!��)	b-��Y%9�Mm[k��u�c���(q��p���vhg>6-�"�?f94]�4>���Ǫ4@�3�B�!�|&#*�Z�m9hÔ��8�˯�@�Yų�E$�\ 
NZ�0/pG�:c�ɮd\H0�,Z�PAG�=�0Y������a��\L"&�m1V$�?�*A�$�̌���7����ܶ�4Qo߽ @�C��2ӗ[������4�����fGiY]N������ 0��Y����f1�%j�x�y�]L�؂�V���QC�L[�BԞE�O58�϶0�'����z[\.J����.N������^��I)��ԋ�3�I5�H>�܍)����Iz�ص�o�SU�}7.h�����r|�LW�w^OM_��Yd����^�]�X����%���t�q8��oŅs��R� ��ѩe���@�)�}�M�g��7Unƾ�&�aL�o[��}��t	e��q�z�޶J�RD�cB!�����F��L�=zp�cfjɬa����f\�yI��$��X.�}Ե<2��cTO�Pl��q9 ؔ!h<D�����.��}�8j��a=ث�R�m��7�̔#��FZ��ṥ���)�S�Pu2�j�8�u�!y�rX��� *�;����)���2�O��
��I/F��{��а��rm^t;~I����KA��mB|?�yg�B΍2\��,��&<ɞ�[HG��� @�f�T+���*gCО��[����5Wy����"�Vκ=��(3�&���y��"�o!�r��kM��c%�h:���.�<�K�.,����&9eȣ�ʯ��?��+�ߠR��.B���`�8�j��w�-=&�ג�?9��E;/��G���iB>㕔���Ԉ4�~k z���0١{*���A^�F�k����,�^6��Fq��K�g���E��#����S%�a���R�?��NƝ��iW,<�:~ *a7b�=ք��)=P���p뗧o���@�����Kd�v,Z�|QĢp�a��
�!!�x,^�μᳰ�GEG�?�i�Օ��ޛq+�%�r�ڄ��	u�y��~�� .>"���^�l�k7�j�Մ����4�k2K����2�_j�e�z��V���Br*�~�eU����9�vt���@��x����qD�K��i��5����؜*�=�
2�I�n/���	r�9�ǵ^S.9�:$�ٶ�+�����]8o��U<|B��:�բN�fQ��5�BZ�}N7e\A��/�y���*y�b7���$��f���bc���d���z��՗H�7��l���N��70\0��z�k�{[c-tN$�������9��eB�F��l�Rɼ?�5�ջ�B��D!lP�#�<p����2y���=�eu�_o�)�G��'��τ~HO������,5�>�]�Ek�Y����g��<�@��8�=eqAt@^6 ӑ�_@#�����b�ί�k��Ö�h�U�!̐ ����ٌ����wp�1�b`lz�a���MksM�!o}Wy�%I����Q�æ�N���$D;�m������J���kP�>l7�8*]�æ�K��}�kO��v�V��\���w#Y�eI���b�����Ϟk- 7��,�l=�g���a������u��~�3��.����-|~Rr&>�;���t�n�Kα .�JO�++q=6$��e+)La
k�3��+ȽCU�SeiC3P�^4��_mO��W�MS���}6�8Ŵ>�q
8dD0�!����;�Ysb��g/Z�#2�L�0�����F�^������.Z�B����{�g��k���
I��~��>
�9+�5�0���5�'f:��5��-o�5}
�3*�C̛z�X�U�_���m��p,����k/h�z&ޱS�҅�M߆'�(��xT~1|C���'�^��5e����cM����P��BduEo�z�R�z� X5�\�j�I^���wxU<�&y����07V'� �vVUE�	�t�i2"�s3�h��A���㚙���]SK�'.��mRW��=��~�,���Z�z����A\���ʆ��[�7Okش�}9 �Io�/h� <pj��d�Ḻ�n���gO���h]78������5q��E?/�kSq\mT���PY�3FKlK�'��a�`%>x��#��&lCրǊLx���C�x�v%zL\c�M[�Rc-\�nU��'Q����Ū�E��KH��* ���驔��ކ�����_5�Ն�0de~&k��*�����Q�����mՊ��%����p~o�N�:m�|ltg�y��[n�}��\Ļ�t yS%ޭW��9�E9�3��p��'�`j�-��l�R=5!S↟���ǜ&�:�����-+B��3 aL<s+O�o�ˊ�wY����T����β�S�#��M��-~eTC���3[�7��'�le������]C��`֩�o�W���ޢ�Ĳi�)LYF"L�o�x�c�?�m3�8�G�Hi�����ǯ���C�)ݠ�e�ڭ'{:�Jˮ�A3�e��;b_��-:ӧKX����E�Q�\�;^����@���ޥ���swb�I���8u[
O�wQ񶱽;�(�	�םer`?��;x���NFO��2:���	����Ie���
F7ZU&ɂ���)���S��`�؁+[1P����9*$����H��n���5־�\��~5�u�!��������}]���eǢU��D�T]Lk7ڙ�1-�BC(Q��E�6����S=�(�T�������omO�g�"����vrn#���AAO/�Z@߉`->�� L�6e���d� 0��U�B:-������[谽�'�@(����'��A�������h	�i�	���]1��W�O�G�9��0E�nӛ)X��L=�݆+����3�V?c9�5ǡP����{�O�8cR	=Rz���3�� d�V풬��<D#�X9�fy���!�`�i2@���KaԮ�ؔ�(�\��%� �����p[/�����5�8�J���E	�-��n��j_>ĕ��`�D2�� ���I0�E�EG�=l�	|��1(��BE#S���k�}�.-RygYI��$� �KMzM�\�'TI���KG=���a'n�޵I����GdDu�2TQ�ӥ�\,	�������S�M	�t�wYc������>��C��Ӊ:�%zN������N�jT�p �&����e���WS�3E�Ml�o��tl�钁"�7o&yU'��jP�m�ٴ�qP~�ƜE�ճ��&��bt��$]֍�1ք�"D���W.�,nZ�UM��>��H�e�T�`��{�^y*EQ�jz�m����&�~�A����i��wQ��r�g���J��]�ϊ	 }����6��w�BL�Z"��&�;�E&�jdd�K��o�P���"���{����M}]D'���ΖC����v)�r�ar���TC�^^�9��+`:ly�7�$��*�t�s�@�&�`�НZ�X��&'Be�[�z��xeR����߭l�{l�尾b���^A�B2��L�DU��� S�'����-�<`����52�sZI�xЎ������j%ʕ�SJ|-ꬑ`&�M�Y�2-#�.�=B��7�"* iK�Տ�[8�++2i,�����I|��&Uǜ�~fZ@�P�'Y|�����/	�-'�;�����1}��j-v�S��7��v<~o���H_h��<��wɖǷχdV1���K�e{�����Ɠ�|-�~!Q���q�[�=6ڥ1?y�&�ʄRg��OU�R���m���h��X�f�&�_�=�"�`T	:�^�4+��PT�g���'�NO�k��xg'W�w�����p���<f�%��N��~ǔ���G�W�D>�H���OP�o�Y��m��� �T� �Y(IB�Z��	k�\��C|H�US)r���B>�����Ľ�\
�g��ם�ԔC�>�k+�G"���[�p��A;�/D����$�;RU\��(�G���Sׅ]����;B���b��L��)%��L]���D.��¤������nB��Z��לH-��+����HoUK�&��a�+�����*�d8��J�_B����ɤʅ�_f����x	ZLB\fF���@ӽ^8o7}a���f�fu���&c��-,��� �'��U���dQ�:eo��<��>k��l�Gw��W�� ���v��@w�W3�sj#;�ҹg��=�"�wh ,�-w2����$N�mc�F��U�Cv���c�C��
��)X7Lj��C�.�*�]�p�n?��}�����=��KO�m-f+�ɑ� `�U�>(0N�P #z�B*��Ip��]�OX�.�s�F�W�੅�Y�[��c��:RD��:`)7ML�x!�(Z�	e!&r脨ܿ�Q��\�]�W�,Џ,��y��=j��5;�������<��9u��$#\l�x�M\�8%�1���zpq%ֆ�6��������md��U�?AYPHng?�o�g,���0Ţd�ĿE��~�֢���$#����?*м�(>b��ifè�:��#2t,��l���)z�C�|������H�gʜ ��e��<�xeO�^�FB�=�_7t�������5�I�qޟbB(���7��`�Ԇ���lF1��H�W �.��K�������&k�v�R��LZ|5O�a�࿸�`H���kz0�X|"��9�#je�w�t`Gn4U�\����� @�Q��*�9Ye�C��y�ƭ��:�n�w�C��{��&����4X�C ⽑�u4ű��B"��o�G��}C���D~q�PQA������#졿���^J��! ���c��jU�Jn�d�҂V�5㝄��s���*:Mp�f-)��z:2��
 -DP��Q�%��2��-����hxo`xu�Y
\e}OKmk�Ѷ��9l���
&/�cj`����	�$��!��rw��	��Ł�%�d6LՓ�,��=E�4�j�Ӽ�	��Pe���`�5���